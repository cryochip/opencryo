magic
tech sky130A
magscale 1 2
timestamp 1624053450
<< nwell >>
rect -1196 -1219 1196 1219
<< pmos >>
rect -1000 -1000 1000 1000
<< pdiff >>
rect -1058 988 -1000 1000
rect -1058 -988 -1046 988
rect -1012 -988 -1000 988
rect -1058 -1000 -1000 -988
rect 1000 988 1058 1000
rect 1000 -988 1012 988
rect 1046 -988 1058 988
rect 1000 -1000 1058 -988
<< pdiffc >>
rect -1046 -988 -1012 988
rect 1012 -988 1046 988
<< nsubdiff >>
rect -1160 1149 -1064 1183
rect 1064 1149 1160 1183
rect -1160 1087 -1126 1149
rect 1126 1087 1160 1149
rect -1160 -1149 -1126 -1087
rect 1126 -1149 1160 -1087
rect -1160 -1183 -1064 -1149
rect 1064 -1183 1160 -1149
<< nsubdiffcont >>
rect -1064 1149 1064 1183
rect -1160 -1087 -1126 1087
rect 1126 -1087 1160 1087
rect -1064 -1183 1064 -1149
<< poly >>
rect -1000 1081 1000 1097
rect -1000 1047 -984 1081
rect 984 1047 1000 1081
rect -1000 1000 1000 1047
rect -1000 -1047 1000 -1000
rect -1000 -1081 -984 -1047
rect 984 -1081 1000 -1047
rect -1000 -1097 1000 -1081
<< polycont >>
rect -984 1047 984 1081
rect -984 -1081 984 -1047
<< locali >>
rect -1160 1149 -1064 1183
rect 1064 1149 1160 1183
rect -1160 1087 -1126 1149
rect 1126 1087 1160 1149
rect -1000 1047 -984 1081
rect 984 1047 1000 1081
rect -1046 988 -1012 1004
rect -1046 -1004 -1012 -988
rect 1012 988 1046 1004
rect 1012 -1004 1046 -988
rect -1000 -1081 -984 -1047
rect 984 -1081 1000 -1047
rect -1160 -1149 -1126 -1087
rect 1126 -1149 1160 -1087
rect -1160 -1183 -1064 -1149
rect 1064 -1183 1160 -1149
<< viali >>
rect -984 1047 984 1081
rect -1046 -988 -1012 988
rect 1012 -988 1046 988
rect -984 -1081 984 -1047
<< metal1 >>
rect -996 1081 996 1087
rect -996 1047 -984 1081
rect 984 1047 996 1081
rect -996 1041 996 1047
rect -1052 988 -1006 1000
rect -1052 -988 -1046 988
rect -1012 -988 -1006 988
rect -1052 -1000 -1006 -988
rect 1006 988 1052 1000
rect 1006 -988 1012 988
rect 1046 -988 1052 988
rect 1006 -1000 1052 -988
rect -996 -1047 996 -1041
rect -996 -1081 -984 -1047
rect 984 -1081 996 -1047
rect -996 -1087 996 -1081
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -1143 -1166 1143 1166
string parameters w 10.0 l 10.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagt 0 viagr 0 viagl 0
string library sky130
<< end >>
