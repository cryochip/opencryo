**.subckt test_nmos G1v8 D1v8 B
*.ipin G1v8
*.ipin D1v8
*.ipin B

.include sky130_nfet_1v8_lvt.mod

Vds D1v8 0 1.8
Vgs G1v8 0 0.8

*XM1 D1v8 G1v8 S 0 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1  nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1

*XM1 D1v8 G1v8 S 0 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1

*M1 D1v8 G1v8 S 0 sky130_fd_pr__nfet_01v8_lvt__model L=0.15 W=1

M1 D1v8 G1v8 S 0 sky130_nfet_1v8_lvt L=0.15 W=10

*XM1 D1v8 G1v8 S 0 skytest 

*.subckt skytest d g s b
*M1 d g s b sky130_nfet_1v8_lvt L=0.15 W=10
*.ends

Vss S 0 0V



.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8_lvt/sky130_fd_pr__nfet_01v8_lvt__tt.pm3.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8_lvt/sky130_fd_pr__nfet_01v8_lvt__tt.corner.spice
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8_lvt/sky130_fd_pr__nfet_01v8_lvt__mismatch.corner.spice
*.include ~/skywater-pdk/libraries/sky130_fd_pr/latest/models/corners/tt.spice

* All models
.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/all.spice

* Corner
*.include ~/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/tt/rf.spice

* this experimental option enables mos model bin
* selection based on W/NF instead of W
.option wnflag=1
.option savecurrents
.control
save all
*@XM1.msky130_fd_pr__nfet_01v8_lvt[gm]
dc vgs 0 1.8 0.001 
*print Vss#branch > output.dat
*write test_nmos.raw

wrdata result.dat Vss#branch
print @M1[gm]

let gm = @M1[gm]

wrdata outN.raw gm



exit

.endc


**** end user architecture code
**.ends
** flattened .save nodes
*.save I(Vss)
.end