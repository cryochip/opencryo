* SPICE3 file created from char.ext - technology: sky130A

.subckt char G BN BP SDN0 SDN1 SDN2 SDN3 SDN4 SDN5 SDN6 SDP0 SDP1 SDP2 SDP3 SDP4 SDP5
+ SDP6
X0 SDP6 G SDP5 BP sky130_fd_pr__pfet_01v8 w=1e+07u l=1e+07u
X1 SDP4 G SDP3 BP sky130_fd_pr__pfet_01v8 w=3e+06u l=600000u
X2 SDN4 G SDN3 BN sky130_fd_pr__nfet_01v8 w=3e+06u l=600000u
X3 SDP5 G SDP4 BP sky130_fd_pr__pfet_01v8 w=3e+06u l=1e+06u
X4 SDN6 G SDN5 BN sky130_fd_pr__nfet_01v8 w=1e+07u l=1e+07u
X5 SDN1 G SDN0 BN sky130_fd_pr__nfet_01v8 w=450000u l=150000u
X6 SDP1 G SDP0 BP sky130_fd_pr__pfet_01v8 w=450000u l=150000u
X7 SDP3 G SDP2 BP sky130_fd_pr__pfet_01v8 w=3e+06u l=300000u
X8 SDP2 G SDP1 BP sky130_fd_pr__pfet_01v8 w=3e+06u l=150000u
X9 SDN2 G SDN1 BN sky130_fd_pr__nfet_01v8 w=3e+06u l=150000u
X10 SDN3 G SDN2 BN sky130_fd_pr__nfet_01v8 w=3e+06u l=300000u
X11 SDN5 G SDN4 BN sky130_fd_pr__nfet_01v8 w=3e+06u l=1e+06u
C0 BP SDP5 2.21fF
.ends

