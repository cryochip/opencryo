magic
tech sky130A
magscale 1 2
timestamp 1624061269
<< pwell >>
rect -1457 -9710 1457 9710
<< nmos >>
rect -1261 -9500 -1061 9500
rect -1003 -9500 -803 9500
rect -745 -9500 -545 9500
rect -487 -9500 -287 9500
rect -229 -9500 -29 9500
rect 29 -9500 229 9500
rect 287 -9500 487 9500
rect 545 -9500 745 9500
rect 803 -9500 1003 9500
rect 1061 -9500 1261 9500
<< ndiff >>
rect -1319 9488 -1261 9500
rect -1319 -9488 -1307 9488
rect -1273 -9488 -1261 9488
rect -1319 -9500 -1261 -9488
rect -1061 9488 -1003 9500
rect -1061 -9488 -1049 9488
rect -1015 -9488 -1003 9488
rect -1061 -9500 -1003 -9488
rect -803 9488 -745 9500
rect -803 -9488 -791 9488
rect -757 -9488 -745 9488
rect -803 -9500 -745 -9488
rect -545 9488 -487 9500
rect -545 -9488 -533 9488
rect -499 -9488 -487 9488
rect -545 -9500 -487 -9488
rect -287 9488 -229 9500
rect -287 -9488 -275 9488
rect -241 -9488 -229 9488
rect -287 -9500 -229 -9488
rect -29 9488 29 9500
rect -29 -9488 -17 9488
rect 17 -9488 29 9488
rect -29 -9500 29 -9488
rect 229 9488 287 9500
rect 229 -9488 241 9488
rect 275 -9488 287 9488
rect 229 -9500 287 -9488
rect 487 9488 545 9500
rect 487 -9488 499 9488
rect 533 -9488 545 9488
rect 487 -9500 545 -9488
rect 745 9488 803 9500
rect 745 -9488 757 9488
rect 791 -9488 803 9488
rect 745 -9500 803 -9488
rect 1003 9488 1061 9500
rect 1003 -9488 1015 9488
rect 1049 -9488 1061 9488
rect 1003 -9500 1061 -9488
rect 1261 9488 1319 9500
rect 1261 -9488 1273 9488
rect 1307 -9488 1319 9488
rect 1261 -9500 1319 -9488
<< ndiffc >>
rect -1307 -9488 -1273 9488
rect -1049 -9488 -1015 9488
rect -791 -9488 -757 9488
rect -533 -9488 -499 9488
rect -275 -9488 -241 9488
rect -17 -9488 17 9488
rect 241 -9488 275 9488
rect 499 -9488 533 9488
rect 757 -9488 791 9488
rect 1015 -9488 1049 9488
rect 1273 -9488 1307 9488
<< psubdiff >>
rect -1421 9640 -1325 9674
rect 1325 9640 1421 9674
rect -1421 9578 -1387 9640
rect 1387 9578 1421 9640
rect -1421 -9640 -1387 -9578
rect 1387 -9640 1421 -9578
rect -1421 -9674 -1325 -9640
rect 1325 -9674 1421 -9640
<< psubdiffcont >>
rect -1325 9640 1325 9674
rect -1421 -9578 -1387 9578
rect 1387 -9578 1421 9578
rect -1325 -9674 1325 -9640
<< poly >>
rect -1261 9572 -1061 9588
rect -1261 9538 -1245 9572
rect -1077 9538 -1061 9572
rect -1261 9500 -1061 9538
rect -1003 9572 -803 9588
rect -1003 9538 -987 9572
rect -819 9538 -803 9572
rect -1003 9500 -803 9538
rect -745 9572 -545 9588
rect -745 9538 -729 9572
rect -561 9538 -545 9572
rect -745 9500 -545 9538
rect -487 9572 -287 9588
rect -487 9538 -471 9572
rect -303 9538 -287 9572
rect -487 9500 -287 9538
rect -229 9572 -29 9588
rect -229 9538 -213 9572
rect -45 9538 -29 9572
rect -229 9500 -29 9538
rect 29 9572 229 9588
rect 29 9538 45 9572
rect 213 9538 229 9572
rect 29 9500 229 9538
rect 287 9572 487 9588
rect 287 9538 303 9572
rect 471 9538 487 9572
rect 287 9500 487 9538
rect 545 9572 745 9588
rect 545 9538 561 9572
rect 729 9538 745 9572
rect 545 9500 745 9538
rect 803 9572 1003 9588
rect 803 9538 819 9572
rect 987 9538 1003 9572
rect 803 9500 1003 9538
rect 1061 9572 1261 9588
rect 1061 9538 1077 9572
rect 1245 9538 1261 9572
rect 1061 9500 1261 9538
rect -1261 -9538 -1061 -9500
rect -1261 -9572 -1245 -9538
rect -1077 -9572 -1061 -9538
rect -1261 -9588 -1061 -9572
rect -1003 -9538 -803 -9500
rect -1003 -9572 -987 -9538
rect -819 -9572 -803 -9538
rect -1003 -9588 -803 -9572
rect -745 -9538 -545 -9500
rect -745 -9572 -729 -9538
rect -561 -9572 -545 -9538
rect -745 -9588 -545 -9572
rect -487 -9538 -287 -9500
rect -487 -9572 -471 -9538
rect -303 -9572 -287 -9538
rect -487 -9588 -287 -9572
rect -229 -9538 -29 -9500
rect -229 -9572 -213 -9538
rect -45 -9572 -29 -9538
rect -229 -9588 -29 -9572
rect 29 -9538 229 -9500
rect 29 -9572 45 -9538
rect 213 -9572 229 -9538
rect 29 -9588 229 -9572
rect 287 -9538 487 -9500
rect 287 -9572 303 -9538
rect 471 -9572 487 -9538
rect 287 -9588 487 -9572
rect 545 -9538 745 -9500
rect 545 -9572 561 -9538
rect 729 -9572 745 -9538
rect 545 -9588 745 -9572
rect 803 -9538 1003 -9500
rect 803 -9572 819 -9538
rect 987 -9572 1003 -9538
rect 803 -9588 1003 -9572
rect 1061 -9538 1261 -9500
rect 1061 -9572 1077 -9538
rect 1245 -9572 1261 -9538
rect 1061 -9588 1261 -9572
<< polycont >>
rect -1245 9538 -1077 9572
rect -987 9538 -819 9572
rect -729 9538 -561 9572
rect -471 9538 -303 9572
rect -213 9538 -45 9572
rect 45 9538 213 9572
rect 303 9538 471 9572
rect 561 9538 729 9572
rect 819 9538 987 9572
rect 1077 9538 1245 9572
rect -1245 -9572 -1077 -9538
rect -987 -9572 -819 -9538
rect -729 -9572 -561 -9538
rect -471 -9572 -303 -9538
rect -213 -9572 -45 -9538
rect 45 -9572 213 -9538
rect 303 -9572 471 -9538
rect 561 -9572 729 -9538
rect 819 -9572 987 -9538
rect 1077 -9572 1245 -9538
<< locali >>
rect -1421 9640 -1325 9674
rect 1325 9640 1421 9674
rect -1421 9578 -1387 9640
rect 1387 9578 1421 9640
rect -1261 9538 -1245 9572
rect -1077 9538 -1061 9572
rect -1003 9538 -987 9572
rect -819 9538 -803 9572
rect -745 9538 -729 9572
rect -561 9538 -545 9572
rect -487 9538 -471 9572
rect -303 9538 -287 9572
rect -229 9538 -213 9572
rect -45 9538 -29 9572
rect 29 9538 45 9572
rect 213 9538 229 9572
rect 287 9538 303 9572
rect 471 9538 487 9572
rect 545 9538 561 9572
rect 729 9538 745 9572
rect 803 9538 819 9572
rect 987 9538 1003 9572
rect 1061 9538 1077 9572
rect 1245 9538 1261 9572
rect -1307 9488 -1273 9504
rect -1307 -9504 -1273 -9488
rect -1049 9488 -1015 9504
rect -1049 -9504 -1015 -9488
rect -791 9488 -757 9504
rect -791 -9504 -757 -9488
rect -533 9488 -499 9504
rect -533 -9504 -499 -9488
rect -275 9488 -241 9504
rect -275 -9504 -241 -9488
rect -17 9488 17 9504
rect -17 -9504 17 -9488
rect 241 9488 275 9504
rect 241 -9504 275 -9488
rect 499 9488 533 9504
rect 499 -9504 533 -9488
rect 757 9488 791 9504
rect 757 -9504 791 -9488
rect 1015 9488 1049 9504
rect 1015 -9504 1049 -9488
rect 1273 9488 1307 9504
rect 1273 -9504 1307 -9488
rect -1261 -9572 -1245 -9538
rect -1077 -9572 -1061 -9538
rect -1003 -9572 -987 -9538
rect -819 -9572 -803 -9538
rect -745 -9572 -729 -9538
rect -561 -9572 -545 -9538
rect -487 -9572 -471 -9538
rect -303 -9572 -287 -9538
rect -229 -9572 -213 -9538
rect -45 -9572 -29 -9538
rect 29 -9572 45 -9538
rect 213 -9572 229 -9538
rect 287 -9572 303 -9538
rect 471 -9572 487 -9538
rect 545 -9572 561 -9538
rect 729 -9572 745 -9538
rect 803 -9572 819 -9538
rect 987 -9572 1003 -9538
rect 1061 -9572 1077 -9538
rect 1245 -9572 1261 -9538
rect -1421 -9640 -1387 -9578
rect 1387 -9640 1421 -9578
rect -1421 -9674 -1325 -9640
rect 1325 -9674 1421 -9640
<< viali >>
rect -1245 9538 -1077 9572
rect -987 9538 -819 9572
rect -729 9538 -561 9572
rect -471 9538 -303 9572
rect -213 9538 -45 9572
rect 45 9538 213 9572
rect 303 9538 471 9572
rect 561 9538 729 9572
rect 819 9538 987 9572
rect 1077 9538 1245 9572
rect -1307 -9488 -1273 9488
rect -1049 -9488 -1015 9488
rect -791 -9488 -757 9488
rect -533 -9488 -499 9488
rect -275 -9488 -241 9488
rect -17 -9488 17 9488
rect 241 -9488 275 9488
rect 499 -9488 533 9488
rect 757 -9488 791 9488
rect 1015 -9488 1049 9488
rect 1273 -9488 1307 9488
rect -1245 -9572 -1077 -9538
rect -987 -9572 -819 -9538
rect -729 -9572 -561 -9538
rect -471 -9572 -303 -9538
rect -213 -9572 -45 -9538
rect 45 -9572 213 -9538
rect 303 -9572 471 -9538
rect 561 -9572 729 -9538
rect 819 -9572 987 -9538
rect 1077 -9572 1245 -9538
<< metal1 >>
rect -1257 9572 -1065 9578
rect -1257 9538 -1245 9572
rect -1077 9538 -1065 9572
rect -1257 9532 -1065 9538
rect -999 9572 -807 9578
rect -999 9538 -987 9572
rect -819 9538 -807 9572
rect -999 9532 -807 9538
rect -741 9572 -549 9578
rect -741 9538 -729 9572
rect -561 9538 -549 9572
rect -741 9532 -549 9538
rect -483 9572 -291 9578
rect -483 9538 -471 9572
rect -303 9538 -291 9572
rect -483 9532 -291 9538
rect -225 9572 -33 9578
rect -225 9538 -213 9572
rect -45 9538 -33 9572
rect -225 9532 -33 9538
rect 33 9572 225 9578
rect 33 9538 45 9572
rect 213 9538 225 9572
rect 33 9532 225 9538
rect 291 9572 483 9578
rect 291 9538 303 9572
rect 471 9538 483 9572
rect 291 9532 483 9538
rect 549 9572 741 9578
rect 549 9538 561 9572
rect 729 9538 741 9572
rect 549 9532 741 9538
rect 807 9572 999 9578
rect 807 9538 819 9572
rect 987 9538 999 9572
rect 807 9532 999 9538
rect 1065 9572 1257 9578
rect 1065 9538 1077 9572
rect 1245 9538 1257 9572
rect 1065 9532 1257 9538
rect -1313 9488 -1267 9500
rect -1313 -9488 -1307 9488
rect -1273 -9488 -1267 9488
rect -1313 -9500 -1267 -9488
rect -1055 9488 -1009 9500
rect -1055 -9488 -1049 9488
rect -1015 -9488 -1009 9488
rect -1055 -9500 -1009 -9488
rect -797 9488 -751 9500
rect -797 -9488 -791 9488
rect -757 -9488 -751 9488
rect -797 -9500 -751 -9488
rect -539 9488 -493 9500
rect -539 -9488 -533 9488
rect -499 -9488 -493 9488
rect -539 -9500 -493 -9488
rect -281 9488 -235 9500
rect -281 -9488 -275 9488
rect -241 -9488 -235 9488
rect -281 -9500 -235 -9488
rect -23 9488 23 9500
rect -23 -9488 -17 9488
rect 17 -9488 23 9488
rect -23 -9500 23 -9488
rect 235 9488 281 9500
rect 235 -9488 241 9488
rect 275 -9488 281 9488
rect 235 -9500 281 -9488
rect 493 9488 539 9500
rect 493 -9488 499 9488
rect 533 -9488 539 9488
rect 493 -9500 539 -9488
rect 751 9488 797 9500
rect 751 -9488 757 9488
rect 791 -9488 797 9488
rect 751 -9500 797 -9488
rect 1009 9488 1055 9500
rect 1009 -9488 1015 9488
rect 1049 -9488 1055 9488
rect 1009 -9500 1055 -9488
rect 1267 9488 1313 9500
rect 1267 -9488 1273 9488
rect 1307 -9488 1313 9488
rect 1267 -9500 1313 -9488
rect -1257 -9538 -1065 -9532
rect -1257 -9572 -1245 -9538
rect -1077 -9572 -1065 -9538
rect -1257 -9578 -1065 -9572
rect -999 -9538 -807 -9532
rect -999 -9572 -987 -9538
rect -819 -9572 -807 -9538
rect -999 -9578 -807 -9572
rect -741 -9538 -549 -9532
rect -741 -9572 -729 -9538
rect -561 -9572 -549 -9538
rect -741 -9578 -549 -9572
rect -483 -9538 -291 -9532
rect -483 -9572 -471 -9538
rect -303 -9572 -291 -9538
rect -483 -9578 -291 -9572
rect -225 -9538 -33 -9532
rect -225 -9572 -213 -9538
rect -45 -9572 -33 -9538
rect -225 -9578 -33 -9572
rect 33 -9538 225 -9532
rect 33 -9572 45 -9538
rect 213 -9572 225 -9538
rect 33 -9578 225 -9572
rect 291 -9538 483 -9532
rect 291 -9572 303 -9538
rect 471 -9572 483 -9538
rect 291 -9578 483 -9572
rect 549 -9538 741 -9532
rect 549 -9572 561 -9538
rect 729 -9572 741 -9538
rect 549 -9578 741 -9572
rect 807 -9538 999 -9532
rect 807 -9572 819 -9538
rect 987 -9572 999 -9538
rect 807 -9578 999 -9572
rect 1065 -9538 1257 -9532
rect 1065 -9572 1077 -9538
rect 1245 -9572 1257 -9538
rect 1065 -9578 1257 -9572
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -1404 -9657 1404 9657
string parameters w 95 l 1 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
