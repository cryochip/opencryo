** VCO Colpitts Oscilator

*.include ~/Circuits/skywater/skywater-pdk/libraries/sky130_fd_pr/latest/models/corners/tt.spice
*.include ~/Circuits/skywater/skywater-pdk/libraries/sky130_fd_pr/latest/models/capacitors/sky130_fd_pr__model__cap_mim.model.spice

.lib "~/Circuits/skywater/skywater-pdk/libraries/sky130_fd_pr/latest/models/sky130.lib.spice" tt

.subckt ColpitOscilator out+ out- *D1v8 G1v8 S1v8 B1v8
*Vosc 5 6 dc 0v sin(0.1 1.0 1k 0) 
*Vran 6 55 trrandom (2 0.5m 0 10m)

*Vosc    5 6  dc 0v sin(0 1.0 5e9)
*VNoi1of 6 55 DC 0 TRNOISE (0 10p 1e-20 12p)

*Vran 6 55 trrandom (2 0.5m 0 10m)

*C1 5 0 0.144p

*XC1 5  0 sky130_fd_pr__cap_mim_m3_2 w=2 l=2 MF=1 *0.144p
*XC2 5  0 sky130_fd_pr__cap_mim_m3_2 w=2 l=2 MF=1 *0.144p
*XC3 5  0 sky130_fd_pr__cap_mim_m3_2 w=4 l=4 MF=1 *0.144p
*XC4 5  0 sky130_fd_pr__cap_mim_m3_2 w=4 l=4 MF=1 *0.144p
*XC5 5  0 sky130_fd_pr__cap_mim_m3_2 w=4 l=4 MF=1 *0.144p

Vdd 1 0 1.8
Vmi out- 0 0

L1  1  55 7n
RL1 55 out+ 73.3

C1 out+ S1v8 0.072p
C2 S1v8 0    0.072p

Vg G1v8 0 1

Ibias S1v8 0 1m

Vb B1v8 0 0

*IIN 5 0 PULSE(0 -0.1 1NS 0.01NS 0.01NS 1NS 100NS)

XM1 out+ G1v8 S1v8 B1v8 sky130_fd_pr__nfet_01v8 L=0.15 W=1.26 ad=W*0.29 pd=2*(W+0.29) as_=W*0.29 ps=2*(W+0.29) nrd=0.29/W nrs=0.29/W sa=0 sb=0 sd=0 nf=1 mult=1
.ends
