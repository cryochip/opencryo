magic
tech sky130A
timestamp 1624076914
<< nwell >>
rect -140 -180 2695 -75
rect 150 -425 2695 -180
rect 1475 -1135 2695 -425
<< nmos >>
rect 0 0 15 45
rect 290 0 305 300
rect 585 0 615 300
rect 895 0 955 300
rect 1235 0 1335 300
rect 1615 0 2615 1000
<< pmos >>
rect 0 -150 15 -105
rect 290 -405 305 -105
rect 585 -405 615 -105
rect 895 -405 955 -105
rect 1235 -405 1335 -105
rect 1615 -1105 2615 -105
<< ndiff >>
rect 1555 955 1615 1000
rect 1555 935 1575 955
rect 1595 935 1615 955
rect 1555 915 1615 935
rect 1555 895 1575 915
rect 1595 895 1615 915
rect 1555 875 1615 895
rect 1555 855 1575 875
rect 1595 855 1615 875
rect 1555 835 1615 855
rect 1555 815 1575 835
rect 1595 815 1615 835
rect 1555 795 1615 815
rect 1555 775 1575 795
rect 1595 775 1615 795
rect 1555 755 1615 775
rect 1555 735 1575 755
rect 1595 735 1615 755
rect 1555 715 1615 735
rect 1555 695 1575 715
rect 1595 695 1615 715
rect 1555 675 1615 695
rect 1555 655 1575 675
rect 1595 655 1615 675
rect 1555 635 1615 655
rect 1555 615 1575 635
rect 1595 615 1615 635
rect 1555 595 1615 615
rect 1555 575 1575 595
rect 1595 575 1615 595
rect 1555 555 1615 575
rect 1555 535 1575 555
rect 1595 535 1615 555
rect 1555 515 1615 535
rect 1555 495 1575 515
rect 1595 495 1615 515
rect 1555 475 1615 495
rect 1555 455 1575 475
rect 1595 455 1615 475
rect 1555 435 1615 455
rect 1555 415 1575 435
rect 1595 415 1615 435
rect 1555 395 1615 415
rect 1555 375 1575 395
rect 1595 375 1615 395
rect 1555 355 1615 375
rect 1555 335 1575 355
rect 1595 335 1615 355
rect 1555 315 1615 335
rect 230 275 290 300
rect 230 255 250 275
rect 270 255 290 275
rect 230 235 290 255
rect 230 215 250 235
rect 270 215 290 235
rect 230 195 290 215
rect 230 175 250 195
rect 270 175 290 195
rect 230 155 290 175
rect 230 135 250 155
rect 270 135 290 155
rect 230 115 290 135
rect 230 95 250 115
rect 270 95 290 115
rect 230 75 290 95
rect 230 55 250 75
rect 270 55 290 75
rect -60 35 0 45
rect -60 15 -40 35
rect -20 15 0 35
rect -60 0 0 15
rect 15 35 75 45
rect 15 15 35 35
rect 55 15 75 35
rect 15 0 75 15
rect 230 35 290 55
rect 230 15 250 35
rect 270 15 290 35
rect 230 0 290 15
rect 305 275 365 300
rect 305 255 325 275
rect 345 255 365 275
rect 305 235 365 255
rect 305 215 325 235
rect 345 215 365 235
rect 305 195 365 215
rect 305 175 325 195
rect 345 175 365 195
rect 305 155 365 175
rect 305 135 325 155
rect 345 135 365 155
rect 305 115 365 135
rect 305 95 325 115
rect 345 95 365 115
rect 305 75 365 95
rect 305 55 325 75
rect 345 55 365 75
rect 305 35 365 55
rect 305 15 325 35
rect 345 15 365 35
rect 305 0 365 15
rect 525 275 585 300
rect 525 255 545 275
rect 565 255 585 275
rect 525 235 585 255
rect 525 215 545 235
rect 565 215 585 235
rect 525 195 585 215
rect 525 175 545 195
rect 565 175 585 195
rect 525 155 585 175
rect 525 135 545 155
rect 565 135 585 155
rect 525 115 585 135
rect 525 95 545 115
rect 565 95 585 115
rect 525 75 585 95
rect 525 55 545 75
rect 565 55 585 75
rect 525 35 585 55
rect 525 15 545 35
rect 565 15 585 35
rect 525 0 585 15
rect 615 275 675 300
rect 615 255 635 275
rect 655 255 675 275
rect 615 235 675 255
rect 615 215 635 235
rect 655 215 675 235
rect 615 195 675 215
rect 615 175 635 195
rect 655 175 675 195
rect 615 155 675 175
rect 615 135 635 155
rect 655 135 675 155
rect 615 115 675 135
rect 615 95 635 115
rect 655 95 675 115
rect 615 75 675 95
rect 615 55 635 75
rect 655 55 675 75
rect 615 35 675 55
rect 615 15 635 35
rect 655 15 675 35
rect 615 0 675 15
rect 835 275 895 300
rect 835 255 855 275
rect 875 255 895 275
rect 835 235 895 255
rect 835 215 855 235
rect 875 215 895 235
rect 835 195 895 215
rect 835 175 855 195
rect 875 175 895 195
rect 835 155 895 175
rect 835 135 855 155
rect 875 135 895 155
rect 835 115 895 135
rect 835 95 855 115
rect 875 95 895 115
rect 835 75 895 95
rect 835 55 855 75
rect 875 55 895 75
rect 835 35 895 55
rect 835 15 855 35
rect 875 15 895 35
rect 835 0 895 15
rect 955 275 1015 300
rect 955 255 975 275
rect 995 255 1015 275
rect 955 235 1015 255
rect 955 215 975 235
rect 995 215 1015 235
rect 955 195 1015 215
rect 955 175 975 195
rect 995 175 1015 195
rect 955 155 1015 175
rect 955 135 975 155
rect 995 135 1015 155
rect 955 115 1015 135
rect 955 95 975 115
rect 995 95 1015 115
rect 955 75 1015 95
rect 955 55 975 75
rect 995 55 1015 75
rect 955 35 1015 55
rect 955 15 975 35
rect 995 15 1015 35
rect 955 0 1015 15
rect 1175 275 1235 300
rect 1175 255 1195 275
rect 1215 255 1235 275
rect 1175 235 1235 255
rect 1175 215 1195 235
rect 1215 215 1235 235
rect 1175 195 1235 215
rect 1175 175 1195 195
rect 1215 175 1235 195
rect 1175 155 1235 175
rect 1175 135 1195 155
rect 1215 135 1235 155
rect 1175 115 1235 135
rect 1175 95 1195 115
rect 1215 95 1235 115
rect 1175 75 1235 95
rect 1175 55 1195 75
rect 1215 55 1235 75
rect 1175 35 1235 55
rect 1175 15 1195 35
rect 1215 15 1235 35
rect 1175 0 1235 15
rect 1335 275 1395 300
rect 1335 255 1355 275
rect 1375 255 1395 275
rect 1335 235 1395 255
rect 1335 215 1355 235
rect 1375 215 1395 235
rect 1335 195 1395 215
rect 1335 175 1355 195
rect 1375 175 1395 195
rect 1335 155 1395 175
rect 1335 135 1355 155
rect 1375 135 1395 155
rect 1335 115 1395 135
rect 1335 95 1355 115
rect 1375 95 1395 115
rect 1335 75 1395 95
rect 1335 55 1355 75
rect 1375 55 1395 75
rect 1335 35 1395 55
rect 1335 15 1355 35
rect 1375 15 1395 35
rect 1335 0 1395 15
rect 1555 295 1575 315
rect 1595 295 1615 315
rect 1555 275 1615 295
rect 1555 255 1575 275
rect 1595 255 1615 275
rect 1555 235 1615 255
rect 1555 215 1575 235
rect 1595 215 1615 235
rect 1555 195 1615 215
rect 1555 175 1575 195
rect 1595 175 1615 195
rect 1555 155 1615 175
rect 1555 135 1575 155
rect 1595 135 1615 155
rect 1555 115 1615 135
rect 1555 95 1575 115
rect 1595 95 1615 115
rect 1555 75 1615 95
rect 1555 55 1575 75
rect 1595 55 1615 75
rect 1555 35 1615 55
rect 1555 15 1575 35
rect 1595 15 1615 35
rect 1555 0 1615 15
rect 2615 955 2675 1000
rect 2615 935 2635 955
rect 2655 935 2675 955
rect 2615 915 2675 935
rect 2615 895 2635 915
rect 2655 895 2675 915
rect 2615 875 2675 895
rect 2615 855 2635 875
rect 2655 855 2675 875
rect 2615 835 2675 855
rect 2615 815 2635 835
rect 2655 815 2675 835
rect 2615 795 2675 815
rect 2615 775 2635 795
rect 2655 775 2675 795
rect 2615 755 2675 775
rect 2615 735 2635 755
rect 2655 735 2675 755
rect 2615 715 2675 735
rect 2615 695 2635 715
rect 2655 695 2675 715
rect 2615 675 2675 695
rect 2615 655 2635 675
rect 2655 655 2675 675
rect 2615 635 2675 655
rect 2615 615 2635 635
rect 2655 615 2675 635
rect 2615 595 2675 615
rect 2615 575 2635 595
rect 2655 575 2675 595
rect 2615 555 2675 575
rect 2615 535 2635 555
rect 2655 535 2675 555
rect 2615 515 2675 535
rect 2615 495 2635 515
rect 2655 495 2675 515
rect 2615 475 2675 495
rect 2615 455 2635 475
rect 2655 455 2675 475
rect 2615 435 2675 455
rect 2615 415 2635 435
rect 2655 415 2675 435
rect 2615 395 2675 415
rect 2615 375 2635 395
rect 2655 375 2675 395
rect 2615 355 2675 375
rect 2615 335 2635 355
rect 2655 335 2675 355
rect 2615 315 2675 335
rect 2615 295 2635 315
rect 2655 295 2675 315
rect 2615 275 2675 295
rect 2615 255 2635 275
rect 2655 255 2675 275
rect 2615 235 2675 255
rect 2615 215 2635 235
rect 2655 215 2675 235
rect 2615 195 2675 215
rect 2615 175 2635 195
rect 2655 175 2675 195
rect 2615 155 2675 175
rect 2615 135 2635 155
rect 2655 135 2675 155
rect 2615 115 2675 135
rect 2615 95 2635 115
rect 2655 95 2675 115
rect 2615 75 2675 95
rect 2615 55 2635 75
rect 2655 55 2675 75
rect 2615 35 2675 55
rect 2615 15 2635 35
rect 2655 15 2675 35
rect 2615 0 2675 15
<< pdiff >>
rect -60 -120 0 -105
rect -60 -140 -40 -120
rect -20 -140 0 -120
rect -60 -150 0 -140
rect 15 -120 75 -105
rect 15 -140 35 -120
rect 55 -140 75 -120
rect 15 -150 75 -140
rect 230 -120 290 -105
rect 230 -140 250 -120
rect 270 -140 290 -120
rect 230 -170 290 -140
rect 230 -190 250 -170
rect 270 -190 290 -170
rect 230 -210 290 -190
rect 230 -230 250 -210
rect 270 -230 290 -210
rect 230 -250 290 -230
rect 230 -270 250 -250
rect 270 -270 290 -250
rect 230 -290 290 -270
rect 230 -310 250 -290
rect 270 -310 290 -290
rect 230 -330 290 -310
rect 230 -350 250 -330
rect 270 -350 290 -330
rect 230 -370 290 -350
rect 230 -390 250 -370
rect 270 -390 290 -370
rect 230 -405 290 -390
rect 305 -120 365 -105
rect 305 -140 325 -120
rect 345 -140 365 -120
rect 305 -170 365 -140
rect 305 -190 325 -170
rect 345 -190 365 -170
rect 305 -210 365 -190
rect 305 -230 325 -210
rect 345 -230 365 -210
rect 305 -250 365 -230
rect 305 -270 325 -250
rect 345 -270 365 -250
rect 305 -290 365 -270
rect 305 -310 325 -290
rect 345 -310 365 -290
rect 305 -330 365 -310
rect 305 -350 325 -330
rect 345 -350 365 -330
rect 305 -370 365 -350
rect 305 -390 325 -370
rect 345 -390 365 -370
rect 305 -405 365 -390
rect 525 -120 585 -105
rect 525 -140 545 -120
rect 565 -140 585 -120
rect 525 -170 585 -140
rect 525 -190 545 -170
rect 565 -190 585 -170
rect 525 -210 585 -190
rect 525 -230 545 -210
rect 565 -230 585 -210
rect 525 -250 585 -230
rect 525 -270 545 -250
rect 565 -270 585 -250
rect 525 -290 585 -270
rect 525 -310 545 -290
rect 565 -310 585 -290
rect 525 -330 585 -310
rect 525 -350 545 -330
rect 565 -350 585 -330
rect 525 -370 585 -350
rect 525 -390 545 -370
rect 565 -390 585 -370
rect 525 -405 585 -390
rect 615 -120 675 -105
rect 615 -140 635 -120
rect 655 -140 675 -120
rect 615 -170 675 -140
rect 615 -190 635 -170
rect 655 -190 675 -170
rect 615 -210 675 -190
rect 615 -230 635 -210
rect 655 -230 675 -210
rect 615 -250 675 -230
rect 615 -270 635 -250
rect 655 -270 675 -250
rect 615 -290 675 -270
rect 615 -310 635 -290
rect 655 -310 675 -290
rect 615 -330 675 -310
rect 615 -350 635 -330
rect 655 -350 675 -330
rect 615 -370 675 -350
rect 615 -390 635 -370
rect 655 -390 675 -370
rect 615 -405 675 -390
rect 835 -120 895 -105
rect 835 -140 855 -120
rect 875 -140 895 -120
rect 835 -170 895 -140
rect 835 -190 855 -170
rect 875 -190 895 -170
rect 835 -210 895 -190
rect 835 -230 855 -210
rect 875 -230 895 -210
rect 835 -250 895 -230
rect 835 -270 855 -250
rect 875 -270 895 -250
rect 835 -290 895 -270
rect 835 -310 855 -290
rect 875 -310 895 -290
rect 835 -330 895 -310
rect 835 -350 855 -330
rect 875 -350 895 -330
rect 835 -370 895 -350
rect 835 -390 855 -370
rect 875 -390 895 -370
rect 835 -405 895 -390
rect 955 -120 1015 -105
rect 955 -140 975 -120
rect 995 -140 1015 -120
rect 955 -170 1015 -140
rect 955 -190 975 -170
rect 995 -190 1015 -170
rect 955 -210 1015 -190
rect 955 -230 975 -210
rect 995 -230 1015 -210
rect 955 -250 1015 -230
rect 955 -270 975 -250
rect 995 -270 1015 -250
rect 955 -290 1015 -270
rect 955 -310 975 -290
rect 995 -310 1015 -290
rect 955 -330 1015 -310
rect 955 -350 975 -330
rect 995 -350 1015 -330
rect 955 -370 1015 -350
rect 955 -390 975 -370
rect 995 -390 1015 -370
rect 955 -405 1015 -390
rect 1175 -120 1235 -105
rect 1175 -140 1195 -120
rect 1215 -140 1235 -120
rect 1175 -170 1235 -140
rect 1175 -190 1195 -170
rect 1215 -190 1235 -170
rect 1175 -210 1235 -190
rect 1175 -230 1195 -210
rect 1215 -230 1235 -210
rect 1175 -250 1235 -230
rect 1175 -270 1195 -250
rect 1215 -270 1235 -250
rect 1175 -290 1235 -270
rect 1175 -310 1195 -290
rect 1215 -310 1235 -290
rect 1175 -330 1235 -310
rect 1175 -350 1195 -330
rect 1215 -350 1235 -330
rect 1175 -370 1235 -350
rect 1175 -390 1195 -370
rect 1215 -390 1235 -370
rect 1175 -405 1235 -390
rect 1335 -120 1395 -105
rect 1335 -140 1355 -120
rect 1375 -140 1395 -120
rect 1335 -170 1395 -140
rect 1335 -190 1355 -170
rect 1375 -190 1395 -170
rect 1335 -210 1395 -190
rect 1335 -230 1355 -210
rect 1375 -230 1395 -210
rect 1335 -250 1395 -230
rect 1335 -270 1355 -250
rect 1375 -270 1395 -250
rect 1335 -290 1395 -270
rect 1335 -310 1355 -290
rect 1375 -310 1395 -290
rect 1335 -330 1395 -310
rect 1335 -350 1355 -330
rect 1375 -350 1395 -330
rect 1335 -370 1395 -350
rect 1335 -390 1355 -370
rect 1375 -390 1395 -370
rect 1335 -405 1395 -390
rect 1555 -120 1615 -105
rect 1555 -140 1575 -120
rect 1595 -140 1615 -120
rect 1555 -190 1615 -140
rect 1555 -210 1575 -190
rect 1595 -210 1615 -190
rect 1555 -230 1615 -210
rect 1555 -250 1575 -230
rect 1595 -250 1615 -230
rect 1555 -270 1615 -250
rect 1555 -290 1575 -270
rect 1595 -290 1615 -270
rect 1555 -310 1615 -290
rect 1555 -330 1575 -310
rect 1595 -330 1615 -310
rect 1555 -350 1615 -330
rect 1555 -370 1575 -350
rect 1595 -370 1615 -350
rect 1555 -390 1615 -370
rect 1555 -410 1575 -390
rect 1595 -410 1615 -390
rect 1555 -430 1615 -410
rect 1555 -450 1575 -430
rect 1595 -450 1615 -430
rect 1555 -470 1615 -450
rect 1555 -490 1575 -470
rect 1595 -490 1615 -470
rect 1555 -510 1615 -490
rect 1555 -530 1575 -510
rect 1595 -530 1615 -510
rect 1555 -550 1615 -530
rect 1555 -570 1575 -550
rect 1595 -570 1615 -550
rect 1555 -590 1615 -570
rect 1555 -610 1575 -590
rect 1595 -610 1615 -590
rect 1555 -630 1615 -610
rect 1555 -650 1575 -630
rect 1595 -650 1615 -630
rect 1555 -670 1615 -650
rect 1555 -690 1575 -670
rect 1595 -690 1615 -670
rect 1555 -710 1615 -690
rect 1555 -730 1575 -710
rect 1595 -730 1615 -710
rect 1555 -750 1615 -730
rect 1555 -770 1575 -750
rect 1595 -770 1615 -750
rect 1555 -790 1615 -770
rect 1555 -810 1575 -790
rect 1595 -810 1615 -790
rect 1555 -830 1615 -810
rect 1555 -850 1575 -830
rect 1595 -850 1615 -830
rect 1555 -870 1615 -850
rect 1555 -890 1575 -870
rect 1595 -890 1615 -870
rect 1555 -910 1615 -890
rect 1555 -930 1575 -910
rect 1595 -930 1615 -910
rect 1555 -950 1615 -930
rect 1555 -970 1575 -950
rect 1595 -970 1615 -950
rect 1555 -990 1615 -970
rect 1555 -1010 1575 -990
rect 1595 -1010 1615 -990
rect 1555 -1030 1615 -1010
rect 1555 -1050 1575 -1030
rect 1595 -1050 1615 -1030
rect 1555 -1070 1615 -1050
rect 1555 -1090 1575 -1070
rect 1595 -1090 1615 -1070
rect 1555 -1105 1615 -1090
rect 2615 -120 2675 -105
rect 2615 -140 2635 -120
rect 2655 -140 2675 -120
rect 2615 -190 2675 -140
rect 2615 -210 2635 -190
rect 2655 -210 2675 -190
rect 2615 -230 2675 -210
rect 2615 -250 2635 -230
rect 2655 -250 2675 -230
rect 2615 -270 2675 -250
rect 2615 -290 2635 -270
rect 2655 -290 2675 -270
rect 2615 -310 2675 -290
rect 2615 -330 2635 -310
rect 2655 -330 2675 -310
rect 2615 -350 2675 -330
rect 2615 -370 2635 -350
rect 2655 -370 2675 -350
rect 2615 -390 2675 -370
rect 2615 -410 2635 -390
rect 2655 -410 2675 -390
rect 2615 -430 2675 -410
rect 2615 -450 2635 -430
rect 2655 -450 2675 -430
rect 2615 -470 2675 -450
rect 2615 -490 2635 -470
rect 2655 -490 2675 -470
rect 2615 -510 2675 -490
rect 2615 -530 2635 -510
rect 2655 -530 2675 -510
rect 2615 -550 2675 -530
rect 2615 -570 2635 -550
rect 2655 -570 2675 -550
rect 2615 -590 2675 -570
rect 2615 -610 2635 -590
rect 2655 -610 2675 -590
rect 2615 -630 2675 -610
rect 2615 -650 2635 -630
rect 2655 -650 2675 -630
rect 2615 -670 2675 -650
rect 2615 -690 2635 -670
rect 2655 -690 2675 -670
rect 2615 -710 2675 -690
rect 2615 -730 2635 -710
rect 2655 -730 2675 -710
rect 2615 -750 2675 -730
rect 2615 -770 2635 -750
rect 2655 -770 2675 -750
rect 2615 -790 2675 -770
rect 2615 -810 2635 -790
rect 2655 -810 2675 -790
rect 2615 -830 2675 -810
rect 2615 -850 2635 -830
rect 2655 -850 2675 -830
rect 2615 -870 2675 -850
rect 2615 -890 2635 -870
rect 2655 -890 2675 -870
rect 2615 -910 2675 -890
rect 2615 -930 2635 -910
rect 2655 -930 2675 -910
rect 2615 -950 2675 -930
rect 2615 -970 2635 -950
rect 2655 -970 2675 -950
rect 2615 -990 2675 -970
rect 2615 -1010 2635 -990
rect 2655 -1010 2675 -990
rect 2615 -1030 2675 -1010
rect 2615 -1050 2635 -1030
rect 2655 -1050 2675 -1030
rect 2615 -1070 2675 -1050
rect 2615 -1090 2635 -1070
rect 2655 -1090 2675 -1070
rect 2615 -1105 2675 -1090
<< ndiffc >>
rect 1575 935 1595 955
rect 1575 895 1595 915
rect 1575 855 1595 875
rect 1575 815 1595 835
rect 1575 775 1595 795
rect 1575 735 1595 755
rect 1575 695 1595 715
rect 1575 655 1595 675
rect 1575 615 1595 635
rect 1575 575 1595 595
rect 1575 535 1595 555
rect 1575 495 1595 515
rect 1575 455 1595 475
rect 1575 415 1595 435
rect 1575 375 1595 395
rect 1575 335 1595 355
rect 250 255 270 275
rect 250 215 270 235
rect 250 175 270 195
rect 250 135 270 155
rect 250 95 270 115
rect 250 55 270 75
rect -40 15 -20 35
rect 35 15 55 35
rect 250 15 270 35
rect 325 255 345 275
rect 325 215 345 235
rect 325 175 345 195
rect 325 135 345 155
rect 325 95 345 115
rect 325 55 345 75
rect 325 15 345 35
rect 545 255 565 275
rect 545 215 565 235
rect 545 175 565 195
rect 545 135 565 155
rect 545 95 565 115
rect 545 55 565 75
rect 545 15 565 35
rect 635 255 655 275
rect 635 215 655 235
rect 635 175 655 195
rect 635 135 655 155
rect 635 95 655 115
rect 635 55 655 75
rect 635 15 655 35
rect 855 255 875 275
rect 855 215 875 235
rect 855 175 875 195
rect 855 135 875 155
rect 855 95 875 115
rect 855 55 875 75
rect 855 15 875 35
rect 975 255 995 275
rect 975 215 995 235
rect 975 175 995 195
rect 975 135 995 155
rect 975 95 995 115
rect 975 55 995 75
rect 975 15 995 35
rect 1195 255 1215 275
rect 1195 215 1215 235
rect 1195 175 1215 195
rect 1195 135 1215 155
rect 1195 95 1215 115
rect 1195 55 1215 75
rect 1195 15 1215 35
rect 1355 255 1375 275
rect 1355 215 1375 235
rect 1355 175 1375 195
rect 1355 135 1375 155
rect 1355 95 1375 115
rect 1355 55 1375 75
rect 1355 15 1375 35
rect 1575 295 1595 315
rect 1575 255 1595 275
rect 1575 215 1595 235
rect 1575 175 1595 195
rect 1575 135 1595 155
rect 1575 95 1595 115
rect 1575 55 1595 75
rect 1575 15 1595 35
rect 2635 935 2655 955
rect 2635 895 2655 915
rect 2635 855 2655 875
rect 2635 815 2655 835
rect 2635 775 2655 795
rect 2635 735 2655 755
rect 2635 695 2655 715
rect 2635 655 2655 675
rect 2635 615 2655 635
rect 2635 575 2655 595
rect 2635 535 2655 555
rect 2635 495 2655 515
rect 2635 455 2655 475
rect 2635 415 2655 435
rect 2635 375 2655 395
rect 2635 335 2655 355
rect 2635 295 2655 315
rect 2635 255 2655 275
rect 2635 215 2655 235
rect 2635 175 2655 195
rect 2635 135 2655 155
rect 2635 95 2655 115
rect 2635 55 2655 75
rect 2635 15 2655 35
<< pdiffc >>
rect -40 -140 -20 -120
rect 35 -140 55 -120
rect 250 -140 270 -120
rect 250 -190 270 -170
rect 250 -230 270 -210
rect 250 -270 270 -250
rect 250 -310 270 -290
rect 250 -350 270 -330
rect 250 -390 270 -370
rect 325 -140 345 -120
rect 325 -190 345 -170
rect 325 -230 345 -210
rect 325 -270 345 -250
rect 325 -310 345 -290
rect 325 -350 345 -330
rect 325 -390 345 -370
rect 545 -140 565 -120
rect 545 -190 565 -170
rect 545 -230 565 -210
rect 545 -270 565 -250
rect 545 -310 565 -290
rect 545 -350 565 -330
rect 545 -390 565 -370
rect 635 -140 655 -120
rect 635 -190 655 -170
rect 635 -230 655 -210
rect 635 -270 655 -250
rect 635 -310 655 -290
rect 635 -350 655 -330
rect 635 -390 655 -370
rect 855 -140 875 -120
rect 855 -190 875 -170
rect 855 -230 875 -210
rect 855 -270 875 -250
rect 855 -310 875 -290
rect 855 -350 875 -330
rect 855 -390 875 -370
rect 975 -140 995 -120
rect 975 -190 995 -170
rect 975 -230 995 -210
rect 975 -270 995 -250
rect 975 -310 995 -290
rect 975 -350 995 -330
rect 975 -390 995 -370
rect 1195 -140 1215 -120
rect 1195 -190 1215 -170
rect 1195 -230 1215 -210
rect 1195 -270 1215 -250
rect 1195 -310 1215 -290
rect 1195 -350 1215 -330
rect 1195 -390 1215 -370
rect 1355 -140 1375 -120
rect 1355 -190 1375 -170
rect 1355 -230 1375 -210
rect 1355 -270 1375 -250
rect 1355 -310 1375 -290
rect 1355 -350 1375 -330
rect 1355 -390 1375 -370
rect 1575 -140 1595 -120
rect 1575 -210 1595 -190
rect 1575 -250 1595 -230
rect 1575 -290 1595 -270
rect 1575 -330 1595 -310
rect 1575 -370 1595 -350
rect 1575 -410 1595 -390
rect 1575 -450 1595 -430
rect 1575 -490 1595 -470
rect 1575 -530 1595 -510
rect 1575 -570 1595 -550
rect 1575 -610 1595 -590
rect 1575 -650 1595 -630
rect 1575 -690 1595 -670
rect 1575 -730 1595 -710
rect 1575 -770 1595 -750
rect 1575 -810 1595 -790
rect 1575 -850 1595 -830
rect 1575 -890 1595 -870
rect 1575 -930 1595 -910
rect 1575 -970 1595 -950
rect 1575 -1010 1595 -990
rect 1575 -1050 1595 -1030
rect 1575 -1090 1595 -1070
rect 2635 -140 2655 -120
rect 2635 -210 2655 -190
rect 2635 -250 2655 -230
rect 2635 -290 2655 -270
rect 2635 -330 2655 -310
rect 2635 -370 2655 -350
rect 2635 -410 2655 -390
rect 2635 -450 2655 -430
rect 2635 -490 2655 -470
rect 2635 -530 2655 -510
rect 2635 -570 2655 -550
rect 2635 -610 2655 -590
rect 2635 -650 2655 -630
rect 2635 -690 2655 -670
rect 2635 -730 2655 -710
rect 2635 -770 2655 -750
rect 2635 -810 2655 -790
rect 2635 -850 2655 -830
rect 2635 -890 2655 -870
rect 2635 -930 2655 -910
rect 2635 -970 2655 -950
rect 2635 -1010 2655 -990
rect 2635 -1050 2655 -1030
rect 2635 -1090 2655 -1070
<< psubdiff >>
rect 1495 955 1555 1000
rect 1495 935 1515 955
rect 1535 935 1555 955
rect 1495 915 1555 935
rect 1495 895 1515 915
rect 1535 895 1555 915
rect 1495 875 1555 895
rect 1495 855 1515 875
rect 1535 855 1555 875
rect 1495 835 1555 855
rect 1495 815 1515 835
rect 1535 815 1555 835
rect 1495 795 1555 815
rect 1495 775 1515 795
rect 1535 775 1555 795
rect 1495 755 1555 775
rect 1495 735 1515 755
rect 1535 735 1555 755
rect 1495 715 1555 735
rect 1495 695 1515 715
rect 1535 695 1555 715
rect 1495 675 1555 695
rect 1495 655 1515 675
rect 1535 655 1555 675
rect 1495 635 1555 655
rect 1495 615 1515 635
rect 1535 615 1555 635
rect 1495 595 1555 615
rect 1495 575 1515 595
rect 1535 575 1555 595
rect 1495 555 1555 575
rect 1495 535 1515 555
rect 1535 535 1555 555
rect 1495 515 1555 535
rect 1495 495 1515 515
rect 1535 495 1555 515
rect 1495 475 1555 495
rect 1495 455 1515 475
rect 1535 455 1555 475
rect 1495 435 1555 455
rect 1495 415 1515 435
rect 1535 415 1555 435
rect 1495 395 1555 415
rect 1495 375 1515 395
rect 1535 375 1555 395
rect 1495 355 1555 375
rect 1495 335 1515 355
rect 1535 335 1555 355
rect 1495 315 1555 335
rect 170 275 230 300
rect 170 255 190 275
rect 210 255 230 275
rect 170 235 230 255
rect 170 215 190 235
rect 210 215 230 235
rect 170 195 230 215
rect 170 175 190 195
rect 210 175 230 195
rect 170 155 230 175
rect 170 135 190 155
rect 210 135 230 155
rect 170 115 230 135
rect 170 95 190 115
rect 210 95 230 115
rect 170 75 230 95
rect 170 55 190 75
rect 210 55 230 75
rect -120 35 -60 45
rect -120 15 -100 35
rect -80 15 -60 35
rect -120 0 -60 15
rect 170 35 230 55
rect 170 15 190 35
rect 210 15 230 35
rect 170 0 230 15
rect 465 275 525 300
rect 465 255 485 275
rect 505 255 525 275
rect 465 235 525 255
rect 465 215 485 235
rect 505 215 525 235
rect 465 195 525 215
rect 465 175 485 195
rect 505 175 525 195
rect 465 155 525 175
rect 465 135 485 155
rect 505 135 525 155
rect 465 115 525 135
rect 465 95 485 115
rect 505 95 525 115
rect 465 75 525 95
rect 465 55 485 75
rect 505 55 525 75
rect 465 35 525 55
rect 465 15 485 35
rect 505 15 525 35
rect 465 0 525 15
rect 775 275 835 300
rect 775 255 795 275
rect 815 255 835 275
rect 775 235 835 255
rect 775 215 795 235
rect 815 215 835 235
rect 775 195 835 215
rect 775 175 795 195
rect 815 175 835 195
rect 775 155 835 175
rect 775 135 795 155
rect 815 135 835 155
rect 775 115 835 135
rect 775 95 795 115
rect 815 95 835 115
rect 775 75 835 95
rect 775 55 795 75
rect 815 55 835 75
rect 775 35 835 55
rect 775 15 795 35
rect 815 15 835 35
rect 775 0 835 15
rect 1115 275 1175 300
rect 1115 255 1135 275
rect 1155 255 1175 275
rect 1115 235 1175 255
rect 1115 215 1135 235
rect 1155 215 1175 235
rect 1115 195 1175 215
rect 1115 175 1135 195
rect 1155 175 1175 195
rect 1115 155 1175 175
rect 1115 135 1135 155
rect 1155 135 1175 155
rect 1115 115 1175 135
rect 1115 95 1135 115
rect 1155 95 1175 115
rect 1115 75 1175 95
rect 1115 55 1135 75
rect 1155 55 1175 75
rect 1115 35 1175 55
rect 1115 15 1135 35
rect 1155 15 1175 35
rect 1115 0 1175 15
rect 1495 295 1515 315
rect 1535 295 1555 315
rect 1495 275 1555 295
rect 1495 255 1515 275
rect 1535 255 1555 275
rect 1495 235 1555 255
rect 1495 215 1515 235
rect 1535 215 1555 235
rect 1495 195 1555 215
rect 1495 175 1515 195
rect 1535 175 1555 195
rect 1495 155 1555 175
rect 1495 135 1515 155
rect 1535 135 1555 155
rect 1495 115 1555 135
rect 1495 95 1515 115
rect 1535 95 1555 115
rect 1495 75 1555 95
rect 1495 55 1515 75
rect 1535 55 1555 75
rect 1495 35 1555 55
rect 1495 15 1515 35
rect 1535 15 1555 35
rect 1495 0 1555 15
<< nsubdiff >>
rect -120 -120 -60 -105
rect -120 -140 -100 -120
rect -80 -140 -60 -120
rect -120 -150 -60 -140
rect 170 -120 230 -105
rect 170 -140 190 -120
rect 210 -140 230 -120
rect 170 -170 230 -140
rect 170 -190 190 -170
rect 210 -190 230 -170
rect 170 -210 230 -190
rect 170 -230 190 -210
rect 210 -230 230 -210
rect 170 -250 230 -230
rect 170 -270 190 -250
rect 210 -270 230 -250
rect 170 -290 230 -270
rect 170 -310 190 -290
rect 210 -310 230 -290
rect 170 -330 230 -310
rect 170 -350 190 -330
rect 210 -350 230 -330
rect 170 -370 230 -350
rect 170 -390 190 -370
rect 210 -390 230 -370
rect 170 -405 230 -390
rect 465 -120 525 -105
rect 465 -140 485 -120
rect 505 -140 525 -120
rect 465 -170 525 -140
rect 465 -190 485 -170
rect 505 -190 525 -170
rect 465 -210 525 -190
rect 465 -230 485 -210
rect 505 -230 525 -210
rect 465 -250 525 -230
rect 465 -270 485 -250
rect 505 -270 525 -250
rect 465 -290 525 -270
rect 465 -310 485 -290
rect 505 -310 525 -290
rect 465 -330 525 -310
rect 465 -350 485 -330
rect 505 -350 525 -330
rect 465 -370 525 -350
rect 465 -390 485 -370
rect 505 -390 525 -370
rect 465 -405 525 -390
rect 775 -120 835 -105
rect 775 -140 795 -120
rect 815 -140 835 -120
rect 775 -170 835 -140
rect 775 -190 795 -170
rect 815 -190 835 -170
rect 775 -210 835 -190
rect 775 -230 795 -210
rect 815 -230 835 -210
rect 775 -250 835 -230
rect 775 -270 795 -250
rect 815 -270 835 -250
rect 775 -290 835 -270
rect 775 -310 795 -290
rect 815 -310 835 -290
rect 775 -330 835 -310
rect 775 -350 795 -330
rect 815 -350 835 -330
rect 775 -370 835 -350
rect 775 -390 795 -370
rect 815 -390 835 -370
rect 775 -405 835 -390
rect 1115 -120 1175 -105
rect 1115 -140 1135 -120
rect 1155 -140 1175 -120
rect 1115 -170 1175 -140
rect 1115 -190 1135 -170
rect 1155 -190 1175 -170
rect 1115 -210 1175 -190
rect 1115 -230 1135 -210
rect 1155 -230 1175 -210
rect 1115 -250 1175 -230
rect 1115 -270 1135 -250
rect 1155 -270 1175 -250
rect 1115 -290 1175 -270
rect 1115 -310 1135 -290
rect 1155 -310 1175 -290
rect 1115 -330 1175 -310
rect 1115 -350 1135 -330
rect 1155 -350 1175 -330
rect 1115 -370 1175 -350
rect 1115 -390 1135 -370
rect 1155 -390 1175 -370
rect 1115 -405 1175 -390
rect 1495 -120 1555 -105
rect 1495 -140 1515 -120
rect 1535 -140 1555 -120
rect 1495 -190 1555 -140
rect 1495 -210 1515 -190
rect 1535 -210 1555 -190
rect 1495 -230 1555 -210
rect 1495 -250 1515 -230
rect 1535 -250 1555 -230
rect 1495 -270 1555 -250
rect 1495 -290 1515 -270
rect 1535 -290 1555 -270
rect 1495 -310 1555 -290
rect 1495 -330 1515 -310
rect 1535 -330 1555 -310
rect 1495 -350 1555 -330
rect 1495 -370 1515 -350
rect 1535 -370 1555 -350
rect 1495 -390 1555 -370
rect 1495 -410 1515 -390
rect 1535 -410 1555 -390
rect 1495 -430 1555 -410
rect 1495 -450 1515 -430
rect 1535 -450 1555 -430
rect 1495 -470 1555 -450
rect 1495 -490 1515 -470
rect 1535 -490 1555 -470
rect 1495 -510 1555 -490
rect 1495 -530 1515 -510
rect 1535 -530 1555 -510
rect 1495 -550 1555 -530
rect 1495 -570 1515 -550
rect 1535 -570 1555 -550
rect 1495 -590 1555 -570
rect 1495 -610 1515 -590
rect 1535 -610 1555 -590
rect 1495 -630 1555 -610
rect 1495 -650 1515 -630
rect 1535 -650 1555 -630
rect 1495 -670 1555 -650
rect 1495 -690 1515 -670
rect 1535 -690 1555 -670
rect 1495 -710 1555 -690
rect 1495 -730 1515 -710
rect 1535 -730 1555 -710
rect 1495 -750 1555 -730
rect 1495 -770 1515 -750
rect 1535 -770 1555 -750
rect 1495 -790 1555 -770
rect 1495 -810 1515 -790
rect 1535 -810 1555 -790
rect 1495 -830 1555 -810
rect 1495 -850 1515 -830
rect 1535 -850 1555 -830
rect 1495 -870 1555 -850
rect 1495 -890 1515 -870
rect 1535 -890 1555 -870
rect 1495 -910 1555 -890
rect 1495 -930 1515 -910
rect 1535 -930 1555 -910
rect 1495 -950 1555 -930
rect 1495 -970 1515 -950
rect 1535 -970 1555 -950
rect 1495 -990 1555 -970
rect 1495 -1010 1515 -990
rect 1535 -1010 1555 -990
rect 1495 -1030 1555 -1010
rect 1495 -1050 1515 -1030
rect 1535 -1050 1555 -1030
rect 1495 -1070 1555 -1050
rect 1495 -1090 1515 -1070
rect 1535 -1090 1555 -1070
rect 1495 -1105 1555 -1090
<< psubdiffcont >>
rect 1515 935 1535 955
rect 1515 895 1535 915
rect 1515 855 1535 875
rect 1515 815 1535 835
rect 1515 775 1535 795
rect 1515 735 1535 755
rect 1515 695 1535 715
rect 1515 655 1535 675
rect 1515 615 1535 635
rect 1515 575 1535 595
rect 1515 535 1535 555
rect 1515 495 1535 515
rect 1515 455 1535 475
rect 1515 415 1535 435
rect 1515 375 1535 395
rect 1515 335 1535 355
rect 190 255 210 275
rect 190 215 210 235
rect 190 175 210 195
rect 190 135 210 155
rect 190 95 210 115
rect 190 55 210 75
rect -100 15 -80 35
rect 190 15 210 35
rect 485 255 505 275
rect 485 215 505 235
rect 485 175 505 195
rect 485 135 505 155
rect 485 95 505 115
rect 485 55 505 75
rect 485 15 505 35
rect 795 255 815 275
rect 795 215 815 235
rect 795 175 815 195
rect 795 135 815 155
rect 795 95 815 115
rect 795 55 815 75
rect 795 15 815 35
rect 1135 255 1155 275
rect 1135 215 1155 235
rect 1135 175 1155 195
rect 1135 135 1155 155
rect 1135 95 1155 115
rect 1135 55 1155 75
rect 1135 15 1155 35
rect 1515 295 1535 315
rect 1515 255 1535 275
rect 1515 215 1535 235
rect 1515 175 1535 195
rect 1515 135 1535 155
rect 1515 95 1535 115
rect 1515 55 1535 75
rect 1515 15 1535 35
<< nsubdiffcont >>
rect -100 -140 -80 -120
rect 190 -140 210 -120
rect 190 -190 210 -170
rect 190 -230 210 -210
rect 190 -270 210 -250
rect 190 -310 210 -290
rect 190 -350 210 -330
rect 190 -390 210 -370
rect 485 -140 505 -120
rect 485 -190 505 -170
rect 485 -230 505 -210
rect 485 -270 505 -250
rect 485 -310 505 -290
rect 485 -350 505 -330
rect 485 -390 505 -370
rect 795 -140 815 -120
rect 795 -190 815 -170
rect 795 -230 815 -210
rect 795 -270 815 -250
rect 795 -310 815 -290
rect 795 -350 815 -330
rect 795 -390 815 -370
rect 1135 -140 1155 -120
rect 1135 -190 1155 -170
rect 1135 -230 1155 -210
rect 1135 -270 1155 -250
rect 1135 -310 1155 -290
rect 1135 -350 1155 -330
rect 1135 -390 1155 -370
rect 1515 -140 1535 -120
rect 1515 -210 1535 -190
rect 1515 -250 1535 -230
rect 1515 -290 1535 -270
rect 1515 -330 1535 -310
rect 1515 -370 1535 -350
rect 1515 -410 1535 -390
rect 1515 -450 1535 -430
rect 1515 -490 1535 -470
rect 1515 -530 1535 -510
rect 1515 -570 1535 -550
rect 1515 -610 1535 -590
rect 1515 -650 1535 -630
rect 1515 -690 1535 -670
rect 1515 -730 1535 -710
rect 1515 -770 1535 -750
rect 1515 -810 1535 -790
rect 1515 -850 1535 -830
rect 1515 -890 1535 -870
rect 1515 -930 1535 -910
rect 1515 -970 1535 -950
rect 1515 -1010 1535 -990
rect 1515 -1050 1535 -1030
rect 1515 -1090 1535 -1070
<< poly >>
rect 1615 1000 2615 1015
rect 290 300 305 315
rect 585 300 615 315
rect 895 300 955 315
rect 1235 300 1335 315
rect 0 45 15 60
rect 0 -25 15 0
rect 290 -25 305 0
rect 585 -25 615 0
rect -40 -35 15 -25
rect -40 -55 -30 -35
rect -10 -55 15 -35
rect -40 -65 15 -55
rect 250 -35 305 -25
rect 250 -55 260 -35
rect 280 -55 305 -35
rect 250 -65 305 -55
rect 545 -35 615 -25
rect 545 -55 555 -35
rect 575 -55 615 -35
rect 545 -65 615 -55
rect 0 -105 15 -65
rect 290 -105 305 -65
rect 585 -105 615 -65
rect 895 -35 955 0
rect 895 -55 915 -35
rect 935 -55 955 -35
rect 895 -105 955 -55
rect 1235 -35 1335 0
rect 1235 -55 1275 -35
rect 1295 -55 1335 -35
rect 1235 -105 1335 -55
rect 1615 -35 2615 0
rect 1615 -55 1655 -35
rect 1675 -55 1730 -35
rect 1750 -55 1805 -35
rect 1825 -55 1880 -35
rect 1900 -55 1955 -35
rect 1975 -55 2030 -35
rect 2050 -55 2105 -35
rect 2125 -55 2180 -35
rect 2200 -55 2255 -35
rect 2275 -55 2330 -35
rect 2350 -55 2405 -35
rect 2425 -55 2480 -35
rect 2500 -55 2555 -35
rect 2575 -55 2615 -35
rect 1615 -105 2615 -55
rect 0 -165 15 -150
rect 290 -420 305 -405
rect 585 -420 615 -405
rect 895 -420 955 -405
rect 1235 -420 1335 -405
rect 1615 -1120 2615 -1105
<< polycont >>
rect -30 -55 -10 -35
rect 260 -55 280 -35
rect 555 -55 575 -35
rect 915 -55 935 -35
rect 1275 -55 1295 -35
rect 1655 -55 1675 -35
rect 1730 -55 1750 -35
rect 1805 -55 1825 -35
rect 1880 -55 1900 -35
rect 1955 -55 1975 -35
rect 2030 -55 2050 -35
rect 2105 -55 2125 -35
rect 2180 -55 2200 -35
rect 2255 -55 2275 -35
rect 2330 -55 2350 -35
rect 2405 -55 2425 -35
rect 2480 -55 2500 -35
rect 2555 -55 2575 -35
<< locali >>
rect 1345 1125 1385 1135
rect 1345 1105 1355 1125
rect 1375 1105 1385 1125
rect 965 935 1005 945
rect 965 915 975 935
rect 995 915 1005 935
rect 625 745 665 755
rect 625 725 635 745
rect 655 725 665 745
rect 315 555 355 565
rect 315 535 325 555
rect 345 535 355 555
rect 25 365 65 375
rect 25 345 35 365
rect 55 345 65 365
rect -110 35 -70 45
rect -110 15 -100 35
rect -80 15 -70 35
rect -110 5 -70 15
rect -50 35 -10 120
rect -50 15 -40 35
rect -20 15 -10 35
rect -50 5 -10 15
rect 25 35 65 345
rect 240 365 280 375
rect 240 345 250 365
rect 270 345 280 365
rect 25 15 35 35
rect 55 15 65 35
rect 25 5 65 15
rect 180 275 220 295
rect 180 255 190 275
rect 210 255 220 275
rect 180 235 220 255
rect 180 215 190 235
rect 210 215 220 235
rect 180 195 220 215
rect 180 175 190 195
rect 210 175 220 195
rect 180 155 220 175
rect 180 135 190 155
rect 210 135 220 155
rect 180 115 220 135
rect 180 95 190 115
rect 210 95 220 115
rect 180 75 220 95
rect 180 55 190 75
rect 210 55 220 75
rect 180 35 220 55
rect 180 15 190 35
rect 210 15 220 35
rect 180 5 220 15
rect 240 275 280 345
rect 240 255 250 275
rect 270 255 280 275
rect 240 235 280 255
rect 240 215 250 235
rect 270 215 280 235
rect 240 195 280 215
rect 240 175 250 195
rect 270 175 280 195
rect 240 155 280 175
rect 240 135 250 155
rect 270 135 280 155
rect 240 115 280 135
rect 240 95 250 115
rect 270 95 280 115
rect 240 75 280 95
rect 240 55 250 75
rect 270 55 280 75
rect 240 35 280 55
rect 240 15 250 35
rect 270 15 280 35
rect 240 5 280 15
rect 315 275 355 535
rect 535 555 575 565
rect 535 535 545 555
rect 565 535 575 555
rect 315 255 325 275
rect 345 255 355 275
rect 315 235 355 255
rect 315 215 325 235
rect 345 215 355 235
rect 315 195 355 215
rect 315 175 325 195
rect 345 175 355 195
rect 315 155 355 175
rect 315 135 325 155
rect 345 135 355 155
rect 315 115 355 135
rect 315 95 325 115
rect 345 95 355 115
rect 315 75 355 95
rect 315 55 325 75
rect 345 55 355 75
rect 315 35 355 55
rect 315 15 325 35
rect 345 15 355 35
rect 315 5 355 15
rect 475 275 515 295
rect 475 255 485 275
rect 505 255 515 275
rect 475 235 515 255
rect 475 215 485 235
rect 505 215 515 235
rect 475 195 515 215
rect 475 175 485 195
rect 505 175 515 195
rect 475 155 515 175
rect 475 135 485 155
rect 505 135 515 155
rect 475 115 515 135
rect 475 95 485 115
rect 505 95 515 115
rect 475 75 515 95
rect 475 55 485 75
rect 505 55 515 75
rect 475 35 515 55
rect 475 15 485 35
rect 505 15 515 35
rect 475 5 515 15
rect 535 275 575 535
rect 535 255 545 275
rect 565 255 575 275
rect 535 235 575 255
rect 535 215 545 235
rect 565 215 575 235
rect 535 195 575 215
rect 535 175 545 195
rect 565 175 575 195
rect 535 155 575 175
rect 535 135 545 155
rect 565 135 575 155
rect 535 115 575 135
rect 535 95 545 115
rect 565 95 575 115
rect 535 75 575 95
rect 535 55 545 75
rect 565 55 575 75
rect 535 35 575 55
rect 535 15 545 35
rect 565 15 575 35
rect 535 5 575 15
rect 625 275 665 725
rect 845 745 885 755
rect 845 725 855 745
rect 875 725 885 745
rect 625 255 635 275
rect 655 255 665 275
rect 625 235 665 255
rect 625 215 635 235
rect 655 215 665 235
rect 625 195 665 215
rect 625 175 635 195
rect 655 175 665 195
rect 625 155 665 175
rect 625 135 635 155
rect 655 135 665 155
rect 625 115 665 135
rect 625 95 635 115
rect 655 95 665 115
rect 625 75 665 95
rect 625 55 635 75
rect 655 55 665 75
rect 625 35 665 55
rect 625 15 635 35
rect 655 15 665 35
rect 625 5 665 15
rect 785 275 825 295
rect 785 255 795 275
rect 815 255 825 275
rect 785 235 825 255
rect 785 215 795 235
rect 815 215 825 235
rect 785 195 825 215
rect 785 175 795 195
rect 815 175 825 195
rect 785 155 825 175
rect 785 135 795 155
rect 815 135 825 155
rect 785 115 825 135
rect 785 95 795 115
rect 815 95 825 115
rect 785 75 825 95
rect 785 55 795 75
rect 815 55 825 75
rect 785 35 825 55
rect 785 15 795 35
rect 815 15 825 35
rect 785 5 825 15
rect 845 275 885 725
rect 845 255 855 275
rect 875 255 885 275
rect 845 235 885 255
rect 845 215 855 235
rect 875 215 885 235
rect 845 195 885 215
rect 845 175 855 195
rect 875 175 885 195
rect 845 155 885 175
rect 845 135 855 155
rect 875 135 885 155
rect 845 115 885 135
rect 845 95 855 115
rect 875 95 885 115
rect 845 75 885 95
rect 845 55 855 75
rect 875 55 885 75
rect 845 35 885 55
rect 845 15 855 35
rect 875 15 885 35
rect 845 5 885 15
rect 965 275 1005 915
rect 1185 935 1225 945
rect 1185 915 1195 935
rect 1215 915 1225 935
rect 965 255 975 275
rect 995 255 1005 275
rect 965 235 1005 255
rect 965 215 975 235
rect 995 215 1005 235
rect 965 195 1005 215
rect 965 175 975 195
rect 995 175 1005 195
rect 965 155 1005 175
rect 965 135 975 155
rect 995 135 1005 155
rect 965 115 1005 135
rect 965 95 975 115
rect 995 95 1005 115
rect 965 75 1005 95
rect 965 55 975 75
rect 995 55 1005 75
rect 965 35 1005 55
rect 965 15 975 35
rect 995 15 1005 35
rect 965 5 1005 15
rect 1125 275 1165 295
rect 1125 255 1135 275
rect 1155 255 1165 275
rect 1125 235 1165 255
rect 1125 215 1135 235
rect 1155 215 1165 235
rect 1125 195 1165 215
rect 1125 175 1135 195
rect 1155 175 1165 195
rect 1125 155 1165 175
rect 1125 135 1135 155
rect 1155 135 1165 155
rect 1125 115 1165 135
rect 1125 95 1135 115
rect 1155 95 1165 115
rect 1125 75 1165 95
rect 1125 55 1135 75
rect 1155 55 1165 75
rect 1125 35 1165 55
rect 1125 15 1135 35
rect 1155 15 1165 35
rect 1125 5 1165 15
rect 1185 275 1225 915
rect 1185 255 1195 275
rect 1215 255 1225 275
rect 1185 235 1225 255
rect 1185 215 1195 235
rect 1215 215 1225 235
rect 1185 195 1225 215
rect 1185 175 1195 195
rect 1215 175 1225 195
rect 1185 155 1225 175
rect 1185 135 1195 155
rect 1215 135 1225 155
rect 1185 115 1225 135
rect 1185 95 1195 115
rect 1215 95 1225 115
rect 1185 75 1225 95
rect 1185 55 1195 75
rect 1215 55 1225 75
rect 1185 35 1225 55
rect 1185 15 1195 35
rect 1215 15 1225 35
rect 1185 5 1225 15
rect 1345 275 1385 1105
rect 1565 1125 1605 1135
rect 1565 1105 1575 1125
rect 1595 1105 1605 1125
rect 1345 255 1355 275
rect 1375 255 1385 275
rect 1345 235 1385 255
rect 1345 215 1355 235
rect 1375 215 1385 235
rect 1345 195 1385 215
rect 1345 175 1355 195
rect 1375 175 1385 195
rect 1345 155 1385 175
rect 1345 135 1355 155
rect 1375 135 1385 155
rect 1345 115 1385 135
rect 1345 95 1355 115
rect 1375 95 1385 115
rect 1345 75 1385 95
rect 1345 55 1355 75
rect 1375 55 1385 75
rect 1345 35 1385 55
rect 1345 15 1355 35
rect 1375 15 1385 35
rect 1345 5 1385 15
rect 1505 955 1545 990
rect 1505 935 1515 955
rect 1535 935 1545 955
rect 1505 915 1545 935
rect 1505 895 1515 915
rect 1535 895 1545 915
rect 1505 875 1545 895
rect 1505 855 1515 875
rect 1535 855 1545 875
rect 1505 835 1545 855
rect 1505 815 1515 835
rect 1535 815 1545 835
rect 1505 795 1545 815
rect 1505 775 1515 795
rect 1535 775 1545 795
rect 1505 755 1545 775
rect 1505 735 1515 755
rect 1535 735 1545 755
rect 1505 715 1545 735
rect 1505 695 1515 715
rect 1535 695 1545 715
rect 1505 675 1545 695
rect 1505 655 1515 675
rect 1535 655 1545 675
rect 1505 635 1545 655
rect 1505 615 1515 635
rect 1535 615 1545 635
rect 1505 595 1545 615
rect 1505 575 1515 595
rect 1535 575 1545 595
rect 1505 555 1545 575
rect 1505 535 1515 555
rect 1535 535 1545 555
rect 1505 515 1545 535
rect 1505 495 1515 515
rect 1535 495 1545 515
rect 1505 475 1545 495
rect 1505 455 1515 475
rect 1535 455 1545 475
rect 1505 435 1545 455
rect 1505 415 1515 435
rect 1535 415 1545 435
rect 1505 395 1545 415
rect 1505 375 1515 395
rect 1535 375 1545 395
rect 1505 355 1545 375
rect 1505 335 1515 355
rect 1535 335 1545 355
rect 1505 315 1545 335
rect 1505 295 1515 315
rect 1535 295 1545 315
rect 1505 275 1545 295
rect 1505 255 1515 275
rect 1535 255 1545 275
rect 1505 235 1545 255
rect 1505 215 1515 235
rect 1535 215 1545 235
rect 1505 195 1545 215
rect 1505 175 1515 195
rect 1535 175 1545 195
rect 1505 155 1545 175
rect 1505 135 1515 155
rect 1535 135 1545 155
rect 1505 115 1545 135
rect 1505 95 1515 115
rect 1535 95 1545 115
rect 1505 75 1545 95
rect 1505 55 1515 75
rect 1535 55 1545 75
rect 1505 35 1545 55
rect 1505 15 1515 35
rect 1535 15 1545 35
rect 1505 5 1545 15
rect 1565 955 1605 1105
rect 1565 935 1575 955
rect 1595 935 1605 955
rect 1565 915 1605 935
rect 1565 895 1575 915
rect 1595 895 1605 915
rect 1565 875 1605 895
rect 1565 855 1575 875
rect 1595 855 1605 875
rect 1565 835 1605 855
rect 1565 815 1575 835
rect 1595 815 1605 835
rect 1565 795 1605 815
rect 1565 775 1575 795
rect 1595 775 1605 795
rect 1565 755 1605 775
rect 1565 735 1575 755
rect 1595 735 1605 755
rect 1565 715 1605 735
rect 1565 695 1575 715
rect 1595 695 1605 715
rect 1565 675 1605 695
rect 1565 655 1575 675
rect 1595 655 1605 675
rect 1565 635 1605 655
rect 1565 615 1575 635
rect 1595 615 1605 635
rect 1565 595 1605 615
rect 1565 575 1575 595
rect 1595 575 1605 595
rect 1565 555 1605 575
rect 1565 535 1575 555
rect 1595 535 1605 555
rect 1565 515 1605 535
rect 1565 495 1575 515
rect 1595 495 1605 515
rect 1565 475 1605 495
rect 1565 455 1575 475
rect 1595 455 1605 475
rect 1565 435 1605 455
rect 1565 415 1575 435
rect 1595 415 1605 435
rect 1565 395 1605 415
rect 1565 375 1575 395
rect 1595 375 1605 395
rect 1565 355 1605 375
rect 1565 335 1575 355
rect 1595 335 1605 355
rect 1565 315 1605 335
rect 1565 295 1575 315
rect 1595 295 1605 315
rect 1565 275 1605 295
rect 1565 255 1575 275
rect 1595 255 1605 275
rect 1565 235 1605 255
rect 1565 215 1575 235
rect 1595 215 1605 235
rect 1565 195 1605 215
rect 1565 175 1575 195
rect 1595 175 1605 195
rect 1565 155 1605 175
rect 1565 135 1575 155
rect 1595 135 1605 155
rect 1565 115 1605 135
rect 1565 95 1575 115
rect 1595 95 1605 115
rect 1565 75 1605 95
rect 1565 55 1575 75
rect 1595 55 1605 75
rect 1565 35 1605 55
rect 1565 15 1575 35
rect 1595 15 1605 35
rect 1565 5 1605 15
rect 2625 955 2665 1135
rect 2625 935 2635 955
rect 2655 935 2665 955
rect 2625 915 2665 935
rect 2625 895 2635 915
rect 2655 895 2665 915
rect 2625 875 2665 895
rect 2625 855 2635 875
rect 2655 855 2665 875
rect 2625 835 2665 855
rect 2625 815 2635 835
rect 2655 815 2665 835
rect 2625 795 2665 815
rect 2625 775 2635 795
rect 2655 775 2665 795
rect 2625 755 2665 775
rect 2625 735 2635 755
rect 2655 735 2665 755
rect 2625 715 2665 735
rect 2625 695 2635 715
rect 2655 695 2665 715
rect 2625 675 2665 695
rect 2625 655 2635 675
rect 2655 655 2665 675
rect 2625 635 2665 655
rect 2625 615 2635 635
rect 2655 615 2665 635
rect 2625 595 2665 615
rect 2625 575 2635 595
rect 2655 575 2665 595
rect 2625 555 2665 575
rect 2625 535 2635 555
rect 2655 535 2665 555
rect 2625 515 2665 535
rect 2625 495 2635 515
rect 2655 495 2665 515
rect 2625 475 2665 495
rect 2625 455 2635 475
rect 2655 455 2665 475
rect 2625 435 2665 455
rect 2625 415 2635 435
rect 2655 415 2665 435
rect 2625 395 2665 415
rect 2625 375 2635 395
rect 2655 375 2665 395
rect 2625 355 2665 375
rect 2625 335 2635 355
rect 2655 335 2665 355
rect 2625 315 2665 335
rect 2625 295 2635 315
rect 2655 295 2665 315
rect 2625 275 2665 295
rect 2625 255 2635 275
rect 2655 255 2665 275
rect 2625 235 2665 255
rect 2625 215 2635 235
rect 2655 215 2665 235
rect 2625 195 2665 215
rect 2625 175 2635 195
rect 2655 175 2665 195
rect 2625 155 2665 175
rect 2625 135 2635 155
rect 2655 135 2665 155
rect 2625 115 2665 135
rect 2625 95 2635 115
rect 2655 95 2665 115
rect 2625 75 2665 95
rect 2625 55 2635 75
rect 2655 55 2665 75
rect 2625 35 2665 55
rect 2625 15 2635 35
rect 2655 15 2665 35
rect 2625 5 2665 15
rect -40 -35 2585 -25
rect -40 -55 -30 -35
rect -10 -55 260 -35
rect 280 -55 555 -35
rect 575 -55 915 -35
rect 935 -55 1275 -35
rect 1295 -55 1655 -35
rect 1675 -55 1730 -35
rect 1750 -55 1805 -35
rect 1825 -55 1880 -35
rect 1900 -55 1955 -35
rect 1975 -55 2030 -35
rect 2050 -55 2105 -35
rect 2125 -55 2180 -35
rect 2200 -55 2255 -35
rect 2275 -55 2330 -35
rect 2350 -55 2405 -35
rect 2425 -55 2480 -35
rect 2500 -55 2555 -35
rect 2575 -55 2585 -35
rect -40 -65 2585 -55
rect -110 -120 -70 -110
rect -110 -140 -100 -120
rect -80 -140 -70 -120
rect -110 -150 -70 -140
rect -50 -120 -10 -110
rect -50 -140 -40 -120
rect -20 -140 -10 -120
rect -50 -225 -10 -140
rect 25 -120 65 -110
rect 25 -140 35 -120
rect 55 -140 65 -120
rect 25 -450 65 -140
rect 180 -120 220 -110
rect 180 -140 190 -120
rect 210 -140 220 -120
rect 180 -170 220 -140
rect 180 -190 190 -170
rect 210 -190 220 -170
rect 180 -210 220 -190
rect 180 -230 190 -210
rect 210 -230 220 -210
rect 180 -250 220 -230
rect 180 -270 190 -250
rect 210 -270 220 -250
rect 180 -290 220 -270
rect 180 -310 190 -290
rect 210 -310 220 -290
rect 180 -330 220 -310
rect 180 -350 190 -330
rect 210 -350 220 -330
rect 180 -370 220 -350
rect 180 -390 190 -370
rect 210 -390 220 -370
rect 180 -400 220 -390
rect 240 -120 280 -110
rect 240 -140 250 -120
rect 270 -140 280 -120
rect 240 -170 280 -140
rect 240 -190 250 -170
rect 270 -190 280 -170
rect 240 -210 280 -190
rect 240 -230 250 -210
rect 270 -230 280 -210
rect 240 -250 280 -230
rect 240 -270 250 -250
rect 270 -270 280 -250
rect 240 -290 280 -270
rect 240 -310 250 -290
rect 270 -310 280 -290
rect 240 -330 280 -310
rect 240 -350 250 -330
rect 270 -350 280 -330
rect 240 -370 280 -350
rect 240 -390 250 -370
rect 270 -390 280 -370
rect 25 -470 35 -450
rect 55 -470 65 -450
rect 25 -480 65 -470
rect 240 -450 280 -390
rect 240 -470 250 -450
rect 270 -470 280 -450
rect 240 -480 280 -470
rect 315 -120 355 -110
rect 315 -140 325 -120
rect 345 -140 355 -120
rect 315 -170 355 -140
rect 315 -190 325 -170
rect 345 -190 355 -170
rect 315 -210 355 -190
rect 315 -230 325 -210
rect 345 -230 355 -210
rect 315 -250 355 -230
rect 315 -270 325 -250
rect 345 -270 355 -250
rect 315 -290 355 -270
rect 315 -310 325 -290
rect 345 -310 355 -290
rect 315 -330 355 -310
rect 315 -350 325 -330
rect 345 -350 355 -330
rect 315 -370 355 -350
rect 315 -390 325 -370
rect 345 -390 355 -370
rect 315 -640 355 -390
rect 475 -120 515 -110
rect 475 -140 485 -120
rect 505 -140 515 -120
rect 475 -170 515 -140
rect 475 -190 485 -170
rect 505 -190 515 -170
rect 475 -210 515 -190
rect 475 -230 485 -210
rect 505 -230 515 -210
rect 475 -250 515 -230
rect 475 -270 485 -250
rect 505 -270 515 -250
rect 475 -290 515 -270
rect 475 -310 485 -290
rect 505 -310 515 -290
rect 475 -330 515 -310
rect 475 -350 485 -330
rect 505 -350 515 -330
rect 475 -370 515 -350
rect 475 -390 485 -370
rect 505 -390 515 -370
rect 475 -400 515 -390
rect 535 -120 575 -110
rect 535 -140 545 -120
rect 565 -140 575 -120
rect 535 -170 575 -140
rect 535 -190 545 -170
rect 565 -190 575 -170
rect 535 -210 575 -190
rect 535 -230 545 -210
rect 565 -230 575 -210
rect 535 -250 575 -230
rect 535 -270 545 -250
rect 565 -270 575 -250
rect 535 -290 575 -270
rect 535 -310 545 -290
rect 565 -310 575 -290
rect 535 -330 575 -310
rect 535 -350 545 -330
rect 565 -350 575 -330
rect 535 -370 575 -350
rect 535 -390 545 -370
rect 565 -390 575 -370
rect 315 -660 325 -640
rect 345 -660 355 -640
rect 315 -670 355 -660
rect 535 -640 575 -390
rect 535 -660 545 -640
rect 565 -660 575 -640
rect 535 -670 575 -660
rect 625 -120 665 -110
rect 625 -140 635 -120
rect 655 -140 665 -120
rect 625 -170 665 -140
rect 625 -190 635 -170
rect 655 -190 665 -170
rect 625 -210 665 -190
rect 625 -230 635 -210
rect 655 -230 665 -210
rect 625 -250 665 -230
rect 625 -270 635 -250
rect 655 -270 665 -250
rect 625 -290 665 -270
rect 625 -310 635 -290
rect 655 -310 665 -290
rect 625 -330 665 -310
rect 625 -350 635 -330
rect 655 -350 665 -330
rect 625 -370 665 -350
rect 625 -390 635 -370
rect 655 -390 665 -370
rect 625 -830 665 -390
rect 785 -120 825 -110
rect 785 -140 795 -120
rect 815 -140 825 -120
rect 785 -170 825 -140
rect 785 -190 795 -170
rect 815 -190 825 -170
rect 785 -210 825 -190
rect 785 -230 795 -210
rect 815 -230 825 -210
rect 785 -250 825 -230
rect 785 -270 795 -250
rect 815 -270 825 -250
rect 785 -290 825 -270
rect 785 -310 795 -290
rect 815 -310 825 -290
rect 785 -330 825 -310
rect 785 -350 795 -330
rect 815 -350 825 -330
rect 785 -370 825 -350
rect 785 -390 795 -370
rect 815 -390 825 -370
rect 785 -400 825 -390
rect 845 -120 885 -110
rect 845 -140 855 -120
rect 875 -140 885 -120
rect 845 -170 885 -140
rect 845 -190 855 -170
rect 875 -190 885 -170
rect 845 -210 885 -190
rect 845 -230 855 -210
rect 875 -230 885 -210
rect 845 -250 885 -230
rect 845 -270 855 -250
rect 875 -270 885 -250
rect 845 -290 885 -270
rect 845 -310 855 -290
rect 875 -310 885 -290
rect 845 -330 885 -310
rect 845 -350 855 -330
rect 875 -350 885 -330
rect 845 -370 885 -350
rect 845 -390 855 -370
rect 875 -390 885 -370
rect 625 -850 635 -830
rect 655 -850 665 -830
rect 625 -860 665 -850
rect 845 -830 885 -390
rect 845 -850 855 -830
rect 875 -850 885 -830
rect 845 -860 885 -850
rect 965 -120 1005 -110
rect 965 -140 975 -120
rect 995 -140 1005 -120
rect 965 -170 1005 -140
rect 965 -190 975 -170
rect 995 -190 1005 -170
rect 965 -210 1005 -190
rect 965 -230 975 -210
rect 995 -230 1005 -210
rect 965 -250 1005 -230
rect 965 -270 975 -250
rect 995 -270 1005 -250
rect 965 -290 1005 -270
rect 965 -310 975 -290
rect 995 -310 1005 -290
rect 965 -330 1005 -310
rect 965 -350 975 -330
rect 995 -350 1005 -330
rect 965 -370 1005 -350
rect 965 -390 975 -370
rect 995 -390 1005 -370
rect 965 -1020 1005 -390
rect 1125 -120 1165 -110
rect 1125 -140 1135 -120
rect 1155 -140 1165 -120
rect 1125 -170 1165 -140
rect 1125 -190 1135 -170
rect 1155 -190 1165 -170
rect 1125 -210 1165 -190
rect 1125 -230 1135 -210
rect 1155 -230 1165 -210
rect 1125 -250 1165 -230
rect 1125 -270 1135 -250
rect 1155 -270 1165 -250
rect 1125 -290 1165 -270
rect 1125 -310 1135 -290
rect 1155 -310 1165 -290
rect 1125 -330 1165 -310
rect 1125 -350 1135 -330
rect 1155 -350 1165 -330
rect 1125 -370 1165 -350
rect 1125 -390 1135 -370
rect 1155 -390 1165 -370
rect 1125 -400 1165 -390
rect 1185 -120 1225 -110
rect 1185 -140 1195 -120
rect 1215 -140 1225 -120
rect 1185 -170 1225 -140
rect 1185 -190 1195 -170
rect 1215 -190 1225 -170
rect 1185 -210 1225 -190
rect 1185 -230 1195 -210
rect 1215 -230 1225 -210
rect 1185 -250 1225 -230
rect 1185 -270 1195 -250
rect 1215 -270 1225 -250
rect 1185 -290 1225 -270
rect 1185 -310 1195 -290
rect 1215 -310 1225 -290
rect 1185 -330 1225 -310
rect 1185 -350 1195 -330
rect 1215 -350 1225 -330
rect 1185 -370 1225 -350
rect 1185 -390 1195 -370
rect 1215 -390 1225 -370
rect 965 -1040 975 -1020
rect 995 -1040 1005 -1020
rect 965 -1050 1005 -1040
rect 1185 -1020 1225 -390
rect 1185 -1040 1195 -1020
rect 1215 -1040 1225 -1020
rect 1185 -1050 1225 -1040
rect 1345 -120 1385 -110
rect 1345 -140 1355 -120
rect 1375 -140 1385 -120
rect 1345 -170 1385 -140
rect 1345 -190 1355 -170
rect 1375 -190 1385 -170
rect 1345 -210 1385 -190
rect 1345 -230 1355 -210
rect 1375 -230 1385 -210
rect 1345 -250 1385 -230
rect 1345 -270 1355 -250
rect 1375 -270 1385 -250
rect 1345 -290 1385 -270
rect 1345 -310 1355 -290
rect 1375 -310 1385 -290
rect 1345 -330 1385 -310
rect 1345 -350 1355 -330
rect 1375 -350 1385 -330
rect 1345 -370 1385 -350
rect 1345 -390 1355 -370
rect 1375 -390 1385 -370
rect 1345 -1210 1385 -390
rect 1505 -120 1545 -110
rect 1505 -140 1515 -120
rect 1535 -140 1545 -120
rect 1505 -190 1545 -140
rect 1505 -210 1515 -190
rect 1535 -210 1545 -190
rect 1505 -230 1545 -210
rect 1505 -250 1515 -230
rect 1535 -250 1545 -230
rect 1505 -270 1545 -250
rect 1505 -290 1515 -270
rect 1535 -290 1545 -270
rect 1505 -310 1545 -290
rect 1505 -330 1515 -310
rect 1535 -330 1545 -310
rect 1505 -350 1545 -330
rect 1505 -370 1515 -350
rect 1535 -370 1545 -350
rect 1505 -390 1545 -370
rect 1505 -410 1515 -390
rect 1535 -410 1545 -390
rect 1505 -430 1545 -410
rect 1505 -450 1515 -430
rect 1535 -450 1545 -430
rect 1505 -470 1545 -450
rect 1505 -490 1515 -470
rect 1535 -490 1545 -470
rect 1505 -510 1545 -490
rect 1505 -530 1515 -510
rect 1535 -530 1545 -510
rect 1505 -550 1545 -530
rect 1505 -570 1515 -550
rect 1535 -570 1545 -550
rect 1505 -590 1545 -570
rect 1505 -610 1515 -590
rect 1535 -610 1545 -590
rect 1505 -630 1545 -610
rect 1505 -650 1515 -630
rect 1535 -650 1545 -630
rect 1505 -670 1545 -650
rect 1505 -690 1515 -670
rect 1535 -690 1545 -670
rect 1505 -710 1545 -690
rect 1505 -730 1515 -710
rect 1535 -730 1545 -710
rect 1505 -750 1545 -730
rect 1505 -770 1515 -750
rect 1535 -770 1545 -750
rect 1505 -790 1545 -770
rect 1505 -810 1515 -790
rect 1535 -810 1545 -790
rect 1505 -830 1545 -810
rect 1505 -850 1515 -830
rect 1535 -850 1545 -830
rect 1505 -870 1545 -850
rect 1505 -890 1515 -870
rect 1535 -890 1545 -870
rect 1505 -910 1545 -890
rect 1505 -930 1515 -910
rect 1535 -930 1545 -910
rect 1505 -950 1545 -930
rect 1505 -970 1515 -950
rect 1535 -970 1545 -950
rect 1505 -990 1545 -970
rect 1505 -1010 1515 -990
rect 1535 -1010 1545 -990
rect 1505 -1030 1545 -1010
rect 1505 -1050 1515 -1030
rect 1535 -1050 1545 -1030
rect 1505 -1070 1545 -1050
rect 1505 -1090 1515 -1070
rect 1535 -1090 1545 -1070
rect 1505 -1100 1545 -1090
rect 1565 -120 1605 -110
rect 1565 -140 1575 -120
rect 1595 -140 1605 -120
rect 1565 -190 1605 -140
rect 1565 -210 1575 -190
rect 1595 -210 1605 -190
rect 1565 -230 1605 -210
rect 1565 -250 1575 -230
rect 1595 -250 1605 -230
rect 1565 -270 1605 -250
rect 1565 -290 1575 -270
rect 1595 -290 1605 -270
rect 1565 -310 1605 -290
rect 1565 -330 1575 -310
rect 1595 -330 1605 -310
rect 1565 -350 1605 -330
rect 1565 -370 1575 -350
rect 1595 -370 1605 -350
rect 1565 -390 1605 -370
rect 1565 -410 1575 -390
rect 1595 -410 1605 -390
rect 1565 -430 1605 -410
rect 1565 -450 1575 -430
rect 1595 -450 1605 -430
rect 1565 -470 1605 -450
rect 1565 -490 1575 -470
rect 1595 -490 1605 -470
rect 1565 -510 1605 -490
rect 1565 -530 1575 -510
rect 1595 -530 1605 -510
rect 1565 -550 1605 -530
rect 1565 -570 1575 -550
rect 1595 -570 1605 -550
rect 1565 -590 1605 -570
rect 1565 -610 1575 -590
rect 1595 -610 1605 -590
rect 1565 -630 1605 -610
rect 1565 -650 1575 -630
rect 1595 -650 1605 -630
rect 1565 -670 1605 -650
rect 1565 -690 1575 -670
rect 1595 -690 1605 -670
rect 1565 -710 1605 -690
rect 1565 -730 1575 -710
rect 1595 -730 1605 -710
rect 1565 -750 1605 -730
rect 1565 -770 1575 -750
rect 1595 -770 1605 -750
rect 1565 -790 1605 -770
rect 1565 -810 1575 -790
rect 1595 -810 1605 -790
rect 1565 -830 1605 -810
rect 1565 -850 1575 -830
rect 1595 -850 1605 -830
rect 1565 -870 1605 -850
rect 1565 -890 1575 -870
rect 1595 -890 1605 -870
rect 1565 -910 1605 -890
rect 1565 -930 1575 -910
rect 1595 -930 1605 -910
rect 1565 -950 1605 -930
rect 1565 -970 1575 -950
rect 1595 -970 1605 -950
rect 1565 -990 1605 -970
rect 1565 -1010 1575 -990
rect 1595 -1010 1605 -990
rect 1565 -1030 1605 -1010
rect 1565 -1050 1575 -1030
rect 1595 -1050 1605 -1030
rect 1565 -1070 1605 -1050
rect 1565 -1090 1575 -1070
rect 1595 -1090 1605 -1070
rect 1345 -1230 1355 -1210
rect 1375 -1230 1385 -1210
rect 1345 -1240 1385 -1230
rect 1565 -1210 1605 -1090
rect 1565 -1230 1575 -1210
rect 1595 -1230 1605 -1210
rect 1565 -1240 1605 -1230
rect 2625 -120 2665 -110
rect 2625 -140 2635 -120
rect 2655 -140 2665 -120
rect 2625 -190 2665 -140
rect 2625 -210 2635 -190
rect 2655 -210 2665 -190
rect 2625 -230 2665 -210
rect 2625 -250 2635 -230
rect 2655 -250 2665 -230
rect 2625 -270 2665 -250
rect 2625 -290 2635 -270
rect 2655 -290 2665 -270
rect 2625 -310 2665 -290
rect 2625 -330 2635 -310
rect 2655 -330 2665 -310
rect 2625 -350 2665 -330
rect 2625 -370 2635 -350
rect 2655 -370 2665 -350
rect 2625 -390 2665 -370
rect 2625 -410 2635 -390
rect 2655 -410 2665 -390
rect 2625 -430 2665 -410
rect 2625 -450 2635 -430
rect 2655 -450 2665 -430
rect 2625 -470 2665 -450
rect 2625 -490 2635 -470
rect 2655 -490 2665 -470
rect 2625 -510 2665 -490
rect 2625 -530 2635 -510
rect 2655 -530 2665 -510
rect 2625 -550 2665 -530
rect 2625 -570 2635 -550
rect 2655 -570 2665 -550
rect 2625 -590 2665 -570
rect 2625 -610 2635 -590
rect 2655 -610 2665 -590
rect 2625 -630 2665 -610
rect 2625 -650 2635 -630
rect 2655 -650 2665 -630
rect 2625 -670 2665 -650
rect 2625 -690 2635 -670
rect 2655 -690 2665 -670
rect 2625 -710 2665 -690
rect 2625 -730 2635 -710
rect 2655 -730 2665 -710
rect 2625 -750 2665 -730
rect 2625 -770 2635 -750
rect 2655 -770 2665 -750
rect 2625 -790 2665 -770
rect 2625 -810 2635 -790
rect 2655 -810 2665 -790
rect 2625 -830 2665 -810
rect 2625 -850 2635 -830
rect 2655 -850 2665 -830
rect 2625 -870 2665 -850
rect 2625 -890 2635 -870
rect 2655 -890 2665 -870
rect 2625 -910 2665 -890
rect 2625 -930 2635 -910
rect 2655 -930 2665 -910
rect 2625 -950 2665 -930
rect 2625 -970 2635 -950
rect 2655 -970 2665 -950
rect 2625 -990 2665 -970
rect 2625 -1010 2635 -990
rect 2655 -1010 2665 -990
rect 2625 -1030 2665 -1010
rect 2625 -1050 2635 -1030
rect 2655 -1050 2665 -1030
rect 2625 -1070 2665 -1050
rect 2625 -1090 2635 -1070
rect 2655 -1090 2665 -1070
rect 2625 -1240 2665 -1090
<< viali >>
rect 1355 1105 1375 1125
rect 975 915 995 935
rect 635 725 655 745
rect 325 535 345 555
rect 35 345 55 365
rect -100 15 -80 35
rect 250 345 270 365
rect 190 15 210 35
rect 545 535 565 555
rect 485 15 505 35
rect 855 725 875 745
rect 795 15 815 35
rect 1195 915 1215 935
rect 1135 15 1155 35
rect 1575 1105 1595 1125
rect 1515 15 1535 35
rect -100 -140 -80 -120
rect 190 -140 210 -120
rect 35 -470 55 -450
rect 250 -470 270 -450
rect 485 -140 505 -120
rect 325 -660 345 -640
rect 545 -660 565 -640
rect 795 -140 815 -120
rect 635 -850 655 -830
rect 855 -850 875 -830
rect 1135 -140 1155 -120
rect 975 -1040 995 -1020
rect 1195 -1040 1215 -1020
rect 1515 -140 1535 -120
rect 1355 -1230 1375 -1210
rect 1575 -1230 1595 -1210
<< metal1 >>
rect 1345 1125 1605 1135
rect 1345 1105 1355 1125
rect 1375 1105 1575 1125
rect 1595 1105 1605 1125
rect 1345 1095 1605 1105
rect 965 935 1225 945
rect 965 915 975 935
rect 995 915 1195 935
rect 1215 915 1225 935
rect 965 905 1225 915
rect 625 745 885 755
rect 625 725 635 745
rect 655 725 855 745
rect 875 725 885 745
rect 625 715 885 725
rect 315 555 575 565
rect 315 535 325 555
rect 345 535 545 555
rect 565 535 575 555
rect 315 525 575 535
rect 25 365 280 375
rect 25 345 35 365
rect 55 345 250 365
rect 270 345 280 365
rect 25 335 280 345
rect -120 35 2695 45
rect -120 15 -100 35
rect -80 15 190 35
rect 210 15 485 35
rect 505 15 795 35
rect 815 15 1135 35
rect 1155 15 1515 35
rect 1535 15 2695 35
rect -120 5 2695 15
rect -140 -120 2695 -110
rect -140 -140 -100 -120
rect -80 -140 190 -120
rect 210 -140 485 -120
rect 505 -140 795 -120
rect 815 -140 1135 -120
rect 1155 -140 1515 -120
rect 1535 -140 2695 -120
rect -140 -150 2695 -140
rect 25 -450 280 -440
rect 25 -470 35 -450
rect 55 -470 250 -450
rect 270 -470 280 -450
rect 25 -480 280 -470
rect 315 -640 575 -630
rect 315 -660 325 -640
rect 345 -660 545 -640
rect 565 -660 575 -640
rect 315 -670 575 -660
rect 625 -830 885 -820
rect 625 -850 635 -830
rect 655 -850 855 -830
rect 875 -850 885 -830
rect 625 -860 885 -850
rect 965 -1020 1225 -1010
rect 965 -1040 975 -1020
rect 995 -1040 1195 -1020
rect 1215 -1040 1225 -1020
rect 965 -1050 1225 -1040
rect 1345 -1210 1605 -1200
rect 1345 -1230 1355 -1210
rect 1375 -1230 1575 -1210
rect 1595 -1230 1605 -1210
rect 1345 -1240 1605 -1230
<< labels >>
rlabel locali -40 -45 -40 -45 7 G
port 1 w
rlabel metal1 -120 25 -120 25 7 BN
port 2 w
rlabel metal1 -140 -130 -140 -130 7 BP
port 3 w
rlabel locali -30 120 -30 120 7 SDN0
port 4 w
rlabel metal1 25 355 25 355 7 SDN1
port 5 w
rlabel metal1 315 545 315 545 7 SDN2
port 6 w
rlabel metal1 625 735 625 735 7 SDN3
port 7 w
rlabel metal1 965 925 965 925 7 SDN4
port 8 w
rlabel metal1 1345 1115 1345 1115 7 SDN5
port 9 w
rlabel locali 2645 1135 2645 1135 7 SDN6
port 10 w
rlabel locali -30 -225 -30 -225 7 SDP0
port 11 w
rlabel metal1 25 -460 25 -460 7 SDP1
port 12 w
rlabel metal1 315 -650 315 -650 7 SDP2
port 13 w
rlabel metal1 625 -840 625 -840 7 SDP3
port 14 w
rlabel metal1 965 -1030 965 -1030 7 SDP4
port 15 w
rlabel metal1 1345 -1220 1345 -1220 7 SDP5
port 16 w
rlabel locali 2645 -1240 2645 -1240 7 SDP6
port 17 w
<< end >>
