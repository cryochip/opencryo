** VCO Colpitts Oscilator

.include ~/Circuits/skywater/skywater-pdk/libraries/sky130_fd_pr/latest/models/corners/tt.spice

.subckt ColpitOscilator 5 55 D1v8 G1v8 S1v8 B1v8
Vosc 5 6 dc 0v sin(0.1 1.0 1k 0) 
Vran 6 55 trrandom (2 0.5m 0 10m)

XM1 D1v8 G1v8 S1v8 B1v8 sky130_fd_pr__nfet_01v8 L=0.15 W=1.26 ad=W*0.29 pd=2*(W+0.29) as_=W*0.29 ps=2*(W+0.29) nrd=0.29/W nrs=0.29/W sa=0 sb=0 sd=0 nf=1 mult=1
.ends
