Source common amplifier

.lib "~/Circuits/skywater/skywater-pdk/libraries/sky130_fd_pr/latest/models/sky130.lib.spice" tt

Vdd 1 0 1.8

*RL1 1 out 73.3

RL1 1 out 662

*Cl out 0 1n

XM1 out G1v8 0 0 sky130_fd_pr__nfet_01v8 L=1 W=95

Ibias 1 G1v8 1m

XM2 G1v8 G1v8 ttt 0 sky130_fd_pr__nfet_01v8 L=1 W=95

C11 in G1v8 1

Vin in 0 0V ac 1

Vtes ttt 0 0V

*.op
.ac dec 1 10 10G

.control
run
print all
print @m.xm2.msky130_fd_pr__nfet_01v8[gm]
* = 4.363036e-03
*print

plot mag(V(out))
*exit
.endc
.end