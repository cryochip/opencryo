magic
tech sky130A
magscale 1 2
timestamp 1624053450
<< nwell >>
rect -256 -519 256 519
<< pmos >>
rect -60 -300 60 300
<< pdiff >>
rect -118 288 -60 300
rect -118 -288 -106 288
rect -72 -288 -60 288
rect -118 -300 -60 -288
rect 60 288 118 300
rect 60 -288 72 288
rect 106 -288 118 288
rect 60 -300 118 -288
<< pdiffc >>
rect -106 -288 -72 288
rect 72 -288 106 288
<< nsubdiff >>
rect -220 449 -124 483
rect 124 449 220 483
rect -220 387 -186 449
rect 186 387 220 449
rect -220 -449 -186 -387
rect 186 -449 220 -387
rect -220 -483 -124 -449
rect 124 -483 220 -449
<< nsubdiffcont >>
rect -124 449 124 483
rect -220 -387 -186 387
rect 186 -387 220 387
rect -124 -483 124 -449
<< poly >>
rect -60 381 60 397
rect -60 347 -44 381
rect 44 347 60 381
rect -60 300 60 347
rect -60 -347 60 -300
rect -60 -381 -44 -347
rect 44 -381 60 -347
rect -60 -397 60 -381
<< polycont >>
rect -44 347 44 381
rect -44 -381 44 -347
<< locali >>
rect -220 449 -124 483
rect 124 449 220 483
rect -220 387 -186 449
rect 186 387 220 449
rect -60 347 -44 381
rect 44 347 60 381
rect -106 288 -72 304
rect -106 -304 -72 -288
rect 72 288 106 304
rect 72 -304 106 -288
rect -60 -381 -44 -347
rect 44 -381 60 -347
rect -220 -449 -186 -387
rect 186 -449 220 -387
rect -220 -483 -124 -449
rect 124 -483 220 -449
<< viali >>
rect -44 347 44 381
rect -106 -288 -72 288
rect 72 -288 106 288
rect -44 -381 44 -347
<< metal1 >>
rect -56 381 56 387
rect -56 347 -44 381
rect 44 347 56 381
rect -56 341 56 347
rect -112 288 -66 300
rect -112 -288 -106 288
rect -72 -288 -66 288
rect -112 -300 -66 -288
rect 66 288 112 300
rect 66 -288 72 288
rect 106 -288 112 288
rect 66 -300 112 -288
rect -56 -347 56 -341
rect -56 -381 -44 -347
rect 44 -381 56 -347
rect -56 -387 56 -381
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -203 -466 203 466
string parameters w 3.0 l 0.6 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagt 0 viagr 0 viagl 0
string library sky130
<< end >>
