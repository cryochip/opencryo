magic
tech sky130A
magscale 1 2
timestamp 1624061269
<< pwell >>
rect -1457 -1160 1457 1160
<< nmos >>
rect -1261 -950 -1061 950
rect -1003 -950 -803 950
rect -745 -950 -545 950
rect -487 -950 -287 950
rect -229 -950 -29 950
rect 29 -950 229 950
rect 287 -950 487 950
rect 545 -950 745 950
rect 803 -950 1003 950
rect 1061 -950 1261 950
<< ndiff >>
rect -1319 938 -1261 950
rect -1319 -938 -1307 938
rect -1273 -938 -1261 938
rect -1319 -950 -1261 -938
rect -1061 938 -1003 950
rect -1061 -938 -1049 938
rect -1015 -938 -1003 938
rect -1061 -950 -1003 -938
rect -803 938 -745 950
rect -803 -938 -791 938
rect -757 -938 -745 938
rect -803 -950 -745 -938
rect -545 938 -487 950
rect -545 -938 -533 938
rect -499 -938 -487 938
rect -545 -950 -487 -938
rect -287 938 -229 950
rect -287 -938 -275 938
rect -241 -938 -229 938
rect -287 -950 -229 -938
rect -29 938 29 950
rect -29 -938 -17 938
rect 17 -938 29 938
rect -29 -950 29 -938
rect 229 938 287 950
rect 229 -938 241 938
rect 275 -938 287 938
rect 229 -950 287 -938
rect 487 938 545 950
rect 487 -938 499 938
rect 533 -938 545 938
rect 487 -950 545 -938
rect 745 938 803 950
rect 745 -938 757 938
rect 791 -938 803 938
rect 745 -950 803 -938
rect 1003 938 1061 950
rect 1003 -938 1015 938
rect 1049 -938 1061 938
rect 1003 -950 1061 -938
rect 1261 938 1319 950
rect 1261 -938 1273 938
rect 1307 -938 1319 938
rect 1261 -950 1319 -938
<< ndiffc >>
rect -1307 -938 -1273 938
rect -1049 -938 -1015 938
rect -791 -938 -757 938
rect -533 -938 -499 938
rect -275 -938 -241 938
rect -17 -938 17 938
rect 241 -938 275 938
rect 499 -938 533 938
rect 757 -938 791 938
rect 1015 -938 1049 938
rect 1273 -938 1307 938
<< psubdiff >>
rect -1421 1090 -1325 1124
rect 1325 1090 1421 1124
rect -1421 1028 -1387 1090
rect 1387 1028 1421 1090
rect -1421 -1090 -1387 -1028
rect 1387 -1090 1421 -1028
rect -1421 -1124 -1325 -1090
rect 1325 -1124 1421 -1090
<< psubdiffcont >>
rect -1325 1090 1325 1124
rect -1421 -1028 -1387 1028
rect 1387 -1028 1421 1028
rect -1325 -1124 1325 -1090
<< poly >>
rect -1261 1022 -1061 1038
rect -1261 988 -1245 1022
rect -1077 988 -1061 1022
rect -1261 950 -1061 988
rect -1003 1022 -803 1038
rect -1003 988 -987 1022
rect -819 988 -803 1022
rect -1003 950 -803 988
rect -745 1022 -545 1038
rect -745 988 -729 1022
rect -561 988 -545 1022
rect -745 950 -545 988
rect -487 1022 -287 1038
rect -487 988 -471 1022
rect -303 988 -287 1022
rect -487 950 -287 988
rect -229 1022 -29 1038
rect -229 988 -213 1022
rect -45 988 -29 1022
rect -229 950 -29 988
rect 29 1022 229 1038
rect 29 988 45 1022
rect 213 988 229 1022
rect 29 950 229 988
rect 287 1022 487 1038
rect 287 988 303 1022
rect 471 988 487 1022
rect 287 950 487 988
rect 545 1022 745 1038
rect 545 988 561 1022
rect 729 988 745 1022
rect 545 950 745 988
rect 803 1022 1003 1038
rect 803 988 819 1022
rect 987 988 1003 1022
rect 803 950 1003 988
rect 1061 1022 1261 1038
rect 1061 988 1077 1022
rect 1245 988 1261 1022
rect 1061 950 1261 988
rect -1261 -988 -1061 -950
rect -1261 -1022 -1245 -988
rect -1077 -1022 -1061 -988
rect -1261 -1038 -1061 -1022
rect -1003 -988 -803 -950
rect -1003 -1022 -987 -988
rect -819 -1022 -803 -988
rect -1003 -1038 -803 -1022
rect -745 -988 -545 -950
rect -745 -1022 -729 -988
rect -561 -1022 -545 -988
rect -745 -1038 -545 -1022
rect -487 -988 -287 -950
rect -487 -1022 -471 -988
rect -303 -1022 -287 -988
rect -487 -1038 -287 -1022
rect -229 -988 -29 -950
rect -229 -1022 -213 -988
rect -45 -1022 -29 -988
rect -229 -1038 -29 -1022
rect 29 -988 229 -950
rect 29 -1022 45 -988
rect 213 -1022 229 -988
rect 29 -1038 229 -1022
rect 287 -988 487 -950
rect 287 -1022 303 -988
rect 471 -1022 487 -988
rect 287 -1038 487 -1022
rect 545 -988 745 -950
rect 545 -1022 561 -988
rect 729 -1022 745 -988
rect 545 -1038 745 -1022
rect 803 -988 1003 -950
rect 803 -1022 819 -988
rect 987 -1022 1003 -988
rect 803 -1038 1003 -1022
rect 1061 -988 1261 -950
rect 1061 -1022 1077 -988
rect 1245 -1022 1261 -988
rect 1061 -1038 1261 -1022
<< polycont >>
rect -1245 988 -1077 1022
rect -987 988 -819 1022
rect -729 988 -561 1022
rect -471 988 -303 1022
rect -213 988 -45 1022
rect 45 988 213 1022
rect 303 988 471 1022
rect 561 988 729 1022
rect 819 988 987 1022
rect 1077 988 1245 1022
rect -1245 -1022 -1077 -988
rect -987 -1022 -819 -988
rect -729 -1022 -561 -988
rect -471 -1022 -303 -988
rect -213 -1022 -45 -988
rect 45 -1022 213 -988
rect 303 -1022 471 -988
rect 561 -1022 729 -988
rect 819 -1022 987 -988
rect 1077 -1022 1245 -988
<< locali >>
rect -1421 1090 -1325 1124
rect 1325 1090 1421 1124
rect -1421 1028 -1387 1090
rect 1387 1028 1421 1090
rect -1261 988 -1245 1022
rect -1077 988 -1061 1022
rect -1003 988 -987 1022
rect -819 988 -803 1022
rect -745 988 -729 1022
rect -561 988 -545 1022
rect -487 988 -471 1022
rect -303 988 -287 1022
rect -229 988 -213 1022
rect -45 988 -29 1022
rect 29 988 45 1022
rect 213 988 229 1022
rect 287 988 303 1022
rect 471 988 487 1022
rect 545 988 561 1022
rect 729 988 745 1022
rect 803 988 819 1022
rect 987 988 1003 1022
rect 1061 988 1077 1022
rect 1245 988 1261 1022
rect -1307 938 -1273 954
rect -1307 -954 -1273 -938
rect -1049 938 -1015 954
rect -1049 -954 -1015 -938
rect -791 938 -757 954
rect -791 -954 -757 -938
rect -533 938 -499 954
rect -533 -954 -499 -938
rect -275 938 -241 954
rect -275 -954 -241 -938
rect -17 938 17 954
rect -17 -954 17 -938
rect 241 938 275 954
rect 241 -954 275 -938
rect 499 938 533 954
rect 499 -954 533 -938
rect 757 938 791 954
rect 757 -954 791 -938
rect 1015 938 1049 954
rect 1015 -954 1049 -938
rect 1273 938 1307 954
rect 1273 -954 1307 -938
rect -1261 -1022 -1245 -988
rect -1077 -1022 -1061 -988
rect -1003 -1022 -987 -988
rect -819 -1022 -803 -988
rect -745 -1022 -729 -988
rect -561 -1022 -545 -988
rect -487 -1022 -471 -988
rect -303 -1022 -287 -988
rect -229 -1022 -213 -988
rect -45 -1022 -29 -988
rect 29 -1022 45 -988
rect 213 -1022 229 -988
rect 287 -1022 303 -988
rect 471 -1022 487 -988
rect 545 -1022 561 -988
rect 729 -1022 745 -988
rect 803 -1022 819 -988
rect 987 -1022 1003 -988
rect 1061 -1022 1077 -988
rect 1245 -1022 1261 -988
rect -1421 -1090 -1387 -1028
rect 1387 -1090 1421 -1028
rect -1421 -1124 -1325 -1090
rect 1325 -1124 1421 -1090
<< viali >>
rect -1245 988 -1077 1022
rect -987 988 -819 1022
rect -729 988 -561 1022
rect -471 988 -303 1022
rect -213 988 -45 1022
rect 45 988 213 1022
rect 303 988 471 1022
rect 561 988 729 1022
rect 819 988 987 1022
rect 1077 988 1245 1022
rect -1307 -938 -1273 938
rect -1049 -938 -1015 938
rect -791 -938 -757 938
rect -533 -938 -499 938
rect -275 -938 -241 938
rect -17 -938 17 938
rect 241 -938 275 938
rect 499 -938 533 938
rect 757 -938 791 938
rect 1015 -938 1049 938
rect 1273 -938 1307 938
rect -1245 -1022 -1077 -988
rect -987 -1022 -819 -988
rect -729 -1022 -561 -988
rect -471 -1022 -303 -988
rect -213 -1022 -45 -988
rect 45 -1022 213 -988
rect 303 -1022 471 -988
rect 561 -1022 729 -988
rect 819 -1022 987 -988
rect 1077 -1022 1245 -988
<< metal1 >>
rect -1257 1022 -1065 1028
rect -1257 988 -1245 1022
rect -1077 988 -1065 1022
rect -1257 982 -1065 988
rect -999 1022 -807 1028
rect -999 988 -987 1022
rect -819 988 -807 1022
rect -999 982 -807 988
rect -741 1022 -549 1028
rect -741 988 -729 1022
rect -561 988 -549 1022
rect -741 982 -549 988
rect -483 1022 -291 1028
rect -483 988 -471 1022
rect -303 988 -291 1022
rect -483 982 -291 988
rect -225 1022 -33 1028
rect -225 988 -213 1022
rect -45 988 -33 1022
rect -225 982 -33 988
rect 33 1022 225 1028
rect 33 988 45 1022
rect 213 988 225 1022
rect 33 982 225 988
rect 291 1022 483 1028
rect 291 988 303 1022
rect 471 988 483 1022
rect 291 982 483 988
rect 549 1022 741 1028
rect 549 988 561 1022
rect 729 988 741 1022
rect 549 982 741 988
rect 807 1022 999 1028
rect 807 988 819 1022
rect 987 988 999 1022
rect 807 982 999 988
rect 1065 1022 1257 1028
rect 1065 988 1077 1022
rect 1245 988 1257 1022
rect 1065 982 1257 988
rect -1313 938 -1267 950
rect -1313 -938 -1307 938
rect -1273 -938 -1267 938
rect -1313 -950 -1267 -938
rect -1055 938 -1009 950
rect -1055 -938 -1049 938
rect -1015 -938 -1009 938
rect -1055 -950 -1009 -938
rect -797 938 -751 950
rect -797 -938 -791 938
rect -757 -938 -751 938
rect -797 -950 -751 -938
rect -539 938 -493 950
rect -539 -938 -533 938
rect -499 -938 -493 938
rect -539 -950 -493 -938
rect -281 938 -235 950
rect -281 -938 -275 938
rect -241 -938 -235 938
rect -281 -950 -235 -938
rect -23 938 23 950
rect -23 -938 -17 938
rect 17 -938 23 938
rect -23 -950 23 -938
rect 235 938 281 950
rect 235 -938 241 938
rect 275 -938 281 938
rect 235 -950 281 -938
rect 493 938 539 950
rect 493 -938 499 938
rect 533 -938 539 938
rect 493 -950 539 -938
rect 751 938 797 950
rect 751 -938 757 938
rect 791 -938 797 938
rect 751 -950 797 -938
rect 1009 938 1055 950
rect 1009 -938 1015 938
rect 1049 -938 1055 938
rect 1009 -950 1055 -938
rect 1267 938 1313 950
rect 1267 -938 1273 938
rect 1307 -938 1313 938
rect 1267 -950 1313 -938
rect -1257 -988 -1065 -982
rect -1257 -1022 -1245 -988
rect -1077 -1022 -1065 -988
rect -1257 -1028 -1065 -1022
rect -999 -988 -807 -982
rect -999 -1022 -987 -988
rect -819 -1022 -807 -988
rect -999 -1028 -807 -1022
rect -741 -988 -549 -982
rect -741 -1022 -729 -988
rect -561 -1022 -549 -988
rect -741 -1028 -549 -1022
rect -483 -988 -291 -982
rect -483 -1022 -471 -988
rect -303 -1022 -291 -988
rect -483 -1028 -291 -1022
rect -225 -988 -33 -982
rect -225 -1022 -213 -988
rect -45 -1022 -33 -988
rect -225 -1028 -33 -1022
rect 33 -988 225 -982
rect 33 -1022 45 -988
rect 213 -1022 225 -988
rect 33 -1028 225 -1022
rect 291 -988 483 -982
rect 291 -1022 303 -988
rect 471 -1022 483 -988
rect 291 -1028 483 -1022
rect 549 -988 741 -982
rect 549 -1022 561 -988
rect 729 -1022 741 -988
rect 549 -1028 741 -1022
rect 807 -988 999 -982
rect 807 -1022 819 -988
rect 987 -1022 999 -988
rect 807 -1028 999 -1022
rect 1065 -988 1257 -982
rect 1065 -1022 1077 -988
rect 1245 -1022 1257 -988
rect 1065 -1028 1257 -1022
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -1404 -1107 1404 1107
string parameters w 9.5 l 1 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
