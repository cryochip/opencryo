magic
tech sky130A
timestamp 1623957158
<< metal4 >>
rect 9960 13294 13315 13315
rect 9960 12696 12696 13294
rect 13294 12696 13315 13294
rect 9960 12675 13315 12696
<< via4 >>
rect 12696 12696 13294 13294
<< metal5 >>
rect 10600 39960 40600 40600
rect 10600 38922 39562 39562
rect 10600 11239 11239 38922
rect 11637 37884 38524 38524
rect 11637 12277 12277 37884
rect 37884 13315 38524 37884
rect 12675 13294 38524 13315
rect 12675 12696 12696 13294
rect 13294 12696 38524 13294
rect 12675 12675 38524 12696
rect 38922 12277 39562 38922
rect 11637 11637 39562 12277
rect 39960 11239 40600 39960
rect 10600 10600 40600 11239
<< end >>
